module note_to_period #(
    parameter int CLOCK_FREQ = 100_000_000
) (
    input logic [6:0] note,
    output logic [24:0] period
);
always_comb begin
    case (note)
        7'd0: period = CLOCK_FREQ / 8.18; // C-1
        7'd1: period = CLOCK_FREQ / 8.66; // C#/Db-1
        7'd2: period = CLOCK_FREQ / 9.18; // D-1
        7'd3: period = CLOCK_FREQ / 9.72; // D#/Eb-1
        7'd4: period = CLOCK_FREQ / 10.30; // E-1
        7'd5: period = CLOCK_FREQ / 10.91; // F-1
        7'd6: period = CLOCK_FREQ / 11.56; // F#/Gb-1
        7'd7: period = CLOCK_FREQ / 12.25; // G-1
        7'd8: period = CLOCK_FREQ / 12.98; // G#/Ab-1
        7'd9: period = CLOCK_FREQ / 13.75; // A-1
        7'd10: period = CLOCK_FREQ / 14.57; // A#/Bb-1
        7'd11: period = CLOCK_FREQ / 15.43; // B-1
        7'd12: period = CLOCK_FREQ / 16.35; // C0
        7'd13: period = CLOCK_FREQ / 17.32; // C#/Db0
        7'd14: period = CLOCK_FREQ / 18.35; // D0
        7'd15: period = CLOCK_FREQ / 19.45; // D#/Eb0
        7'd16: period = CLOCK_FREQ / 20.60; // E0
        7'd17: period = CLOCK_FREQ / 21.83; // F0
        7'd18: period = CLOCK_FREQ / 23.12; // F#/Gb0
        7'd19: period = CLOCK_FREQ / 24.50; // G0
        7'd20: period = CLOCK_FREQ / 25.96; // G#/Ab0
        7'd21: period = CLOCK_FREQ / 27.50; // A0
        7'd22: period = CLOCK_FREQ / 29.14; // A#/Bb0
        7'd23: period = CLOCK_FREQ / 30.87; // B0
        7'd24: period = CLOCK_FREQ / 32.70; // C1
        7'd25: period = CLOCK_FREQ / 34.65; // C#/Db1
        7'd26: period = CLOCK_FREQ / 36.71; // D1
        7'd27: period = CLOCK_FREQ / 38.89; // D#/Eb1
        7'd28: period = CLOCK_FREQ / 41.20; // E1
        7'd29: period = CLOCK_FREQ / 43.65; // F1
        7'd30: period = CLOCK_FREQ / 46.25; // F#/Gb1
        7'd31: period = CLOCK_FREQ / 49.00; // G1
        7'd32: period = CLOCK_FREQ / 51.91; // G#/Ab1
        7'd33: period = CLOCK_FREQ / 55.00; // A1
        7'd34: period = CLOCK_FREQ / 58.27; // A#/Bb1
        7'd35: period = CLOCK_FREQ / 61.74; // B1
        7'd36: period = CLOCK_FREQ / 65.41; // C2
        7'd37: period = CLOCK_FREQ / 69.30; // C#/Db2
        7'd38: period = CLOCK_FREQ / 73.42; // D2
        7'd39: period = CLOCK_FREQ / 77.78; // D#/Eb2
        7'd40: period = CLOCK_FREQ / 82.41; // E2
        7'd41: period = CLOCK_FREQ / 87.31; // F2
        7'd42: period = CLOCK_FREQ / 92.50; // F#/Gb2
        7'd43: period = CLOCK_FREQ / 98.00; // G2
        7'd44: period = CLOCK_FREQ / 103.83; // G#/Ab2
        7'd45: period = CLOCK_FREQ / 110.00; // A2
        7'd46: period = CLOCK_FREQ / 116.54; // A#/Bb2
        7'd47: period = CLOCK_FREQ / 123.47; // B2
        7'd48: period = CLOCK_FREQ / 130.81; // C3
        7'd49: period = CLOCK_FREQ / 138.59; // C#/Db3
        7'd50: period = CLOCK_FREQ / 146.83; // D3
        7'd51: period = CLOCK_FREQ / 155.56; // D#/Eb3
        7'd52: period = CLOCK_FREQ / 164.81; // E3
        7'd53: period = CLOCK_FREQ / 174.61; // F3
        7'd54: period = CLOCK_FREQ / 185.00; // F#/Gb3
        7'd55: period = CLOCK_FREQ / 196.00; // G3
        7'd56: period = CLOCK_FREQ / 207.65; // G#/Ab3
        7'd57: period = CLOCK_FREQ / 220.00; // A3
        7'd58: period = CLOCK_FREQ / 233.08; // A#/Bb3
        7'd59: period = CLOCK_FREQ / 246.94; // B3
        7'd60: period = CLOCK_FREQ / 261.63; // C4 (Middle C)
        7'd61: period = CLOCK_FREQ / 277.18; // C#/Db4
        7'd62: period = CLOCK_FREQ / 293.66; // D4
        7'd63: period = CLOCK_FREQ / 311.13; // D#/Eb4
        7'd64: period = CLOCK_FREQ / 329.63; // E4
        7'd65: period = CLOCK_FREQ / 349.23; // F4
        7'd66: period = CLOCK_FREQ / 369.99; // F#/Gb4
        7'd67: period = CLOCK_FREQ / 392.00; // G4
        7'd68: period = CLOCK_FREQ / 415.30; // G#/Ab4
        7'd69: period = CLOCK_FREQ / 440.00; // A4 (standard tuning)
        7'd70: period = CLOCK_FREQ / 466.16; // A#/Bb4
        7'd71: period = CLOCK_FREQ / 493.88; // B4
        7'd72: period = CLOCK_FREQ / 523.25; // C5
        7'd73: period = CLOCK_FREQ / 554.37; // C#/Db5
        7'd74: period = CLOCK_FREQ / 587.33; // D5
        7'd75: period = CLOCK_FREQ / 622.25; // D#/Eb5
        7'd76: period = CLOCK_FREQ / 659.25; // E5
        7'd77: period = CLOCK_FREQ / 698.46; // F5
        7'd78: period = CLOCK_FREQ / 739.99; // F#/Gb5
        7'd79: period = CLOCK_FREQ / 783.99; // G5
        7'd80: period = CLOCK_FREQ / 830.61; // G#/Ab5
        7'd81: period = CLOCK_FREQ / 880.00; // A5
        7'd82: period = CLOCK_FREQ / 932.33; // A#/Bb5
        7'd83: period = CLOCK_FREQ / 987.77; // B5
        7'd84: period = CLOCK_FREQ / 1046.50; // C6
        7'd85: period = CLOCK_FREQ / 1108.73; // C#/Db6
        7'd86: period = CLOCK_FREQ / 1174.66; // D6
        7'd87: period = CLOCK_FREQ / 1244.51; // D#/Eb6
        7'd88: period = CLOCK_FREQ / 1318.51; // E6
        7'd89: period = CLOCK_FREQ / 1396.91; // F6
        7'd90: period = CLOCK_FREQ / 1479.98; // F#/Gb6
        7'd91: period = CLOCK_FREQ / 1567.98; // G6
        7'd92: period = CLOCK_FREQ / 1661.22; // G#/Ab6
        7'd93: period = CLOCK_FREQ / 1760.00; // A6
        7'd94: period = CLOCK_FREQ / 1864.66; // A#/Bb6
        7'd95: period = CLOCK_FREQ / 1975.53; // B6
        7'd96: period = CLOCK_FREQ / 2093.00; // C7
        7'd97: period = CLOCK_FREQ / 2217.46; // C#/Db7
        7'd98: period = CLOCK_FREQ / 2349.32; // D7
        7'd99: period = CLOCK_FREQ / 2489.02; // D#/Eb7
        7'd100: period = CLOCK_FREQ / 2637.02; // E7
        7'd101: period = CLOCK_FREQ / 2793.83; // F7
        7'd102: period = CLOCK_FREQ / 2959.96; // F#/Gb7
        7'd103: period = CLOCK_FREQ / 3135.96; // G7
        7'd104: period = CLOCK_FREQ / 3322.44; // G#/Ab7
        7'd105: period = CLOCK_FREQ / 3520.00; // A7
        7'd106: period = CLOCK_FREQ / 3729.31; // A#/Bb7
        7'd107: period = CLOCK_FREQ / 3951.07; // B7
        7'd108: period = CLOCK_FREQ / 4186.01; // C8
        7'd109: period = CLOCK_FREQ / 4434.92; // C#/Db8
        7'd110: period = CLOCK_FREQ / 4698.64; // D8
        7'd111: period = CLOCK_FREQ / 4978.03; // D#/Eb8
        7'd112: period = CLOCK_FREQ / 5274.04; // E8
        7'd113: period = CLOCK_FREQ / 5587.65; // F8
        7'd114: period = CLOCK_FREQ / 5919.91; // F#/Gb8
        7'd115: period = CLOCK_FREQ / 6271.93; // G8
        7'd116: period = CLOCK_FREQ / 6644.88; // G#/Ab8
        7'd117: period = CLOCK_FREQ / 7040.00; // A8
        7'd118: period = CLOCK_FREQ / 7458.62; // A#/Bb8
        7'd119: period = CLOCK_FREQ / 7902.13; // B8
        7'd120: period = CLOCK_FREQ / 8372.02; // C9
        7'd121: period = CLOCK_FREQ / 8869.84; // C#/Db9
        7'd122: period = CLOCK_FREQ / 9397.27; // D9
        7'd123: period = CLOCK_FREQ / 9956.06; // D#/Eb9
        7'd124: period = CLOCK_FREQ / 10548.08; // E9
        7'd125: period = CLOCK_FREQ / 11175.30; // F9
        7'd126: period = CLOCK_FREQ / 11839.82; // F#/Gb9
        7'd127: period = CLOCK_FREQ / 12543.85; // G9
        default: period = 32'h0;
    endcase
end       
endmodule