module song5_dur #(
	parameter int CLOCK_FREQ = 100_000_000
) (
	input logic [10:0] note_index,
	output logic [28:0] note_dur // max 10s at 100MHz clock
);

localparam real TEMPO_BPM = 120;
localparam real CYCLES_PER_BEAT = CLOCK_FREQ*(60/TEMPO_BPM);
localparam real CYCLES_PER_US = CLOCK_FREQ/1000_000;

always_comb begin
	// the quarter note is one beat and therfore can be multipled by CYCLES_PER_BEAT
	case (note_index)
		0: note_dur = CYCLES_PER_US * 186719;
		1: note_dur = CYCLES_PER_US * 781;
		2: note_dur = CYCLES_PER_US * 186719;
		3: note_dur = CYCLES_PER_US * 781;
		4: note_dur = CYCLES_PER_US * 186719;
		5: note_dur = CYCLES_PER_US * 781;
		6: note_dur = CYCLES_PER_US * 186719;
		7: note_dur = CYCLES_PER_US * 781;
		8: note_dur = CYCLES_PER_US * 186719;
		9: note_dur = CYCLES_PER_US * 781;
		10: note_dur = CYCLES_PER_US * 186719;
		11: note_dur = CYCLES_PER_US * 781;
		12: note_dur = CYCLES_PER_US * 186719;
		13: note_dur = CYCLES_PER_US * 781;
		14: note_dur = CYCLES_PER_US * 186719;
		15: note_dur = CYCLES_PER_US * 781;
		16: note_dur = CYCLES_PER_US * 374219;
		17: note_dur = CYCLES_PER_US * 781;
		18: note_dur = CYCLES_PER_US * 186719;
		19: note_dur = CYCLES_PER_US * 781;
		20: note_dur = CYCLES_PER_US * 92969;
		21: note_dur = CYCLES_PER_US * 781;
		22: note_dur = CYCLES_PER_US * 92969;
		23: note_dur = CYCLES_PER_US * 781;
		24: note_dur = CYCLES_PER_US * 374219;
		25: note_dur = CYCLES_PER_US * 781;
		26: note_dur = CYCLES_PER_US * 1124219;
		27: note_dur = CYCLES_PER_US * 781;
		28: note_dur = CYCLES_PER_US * 92969;
		29: note_dur = CYCLES_PER_US * 781;
		30: note_dur = CYCLES_PER_US * 92969;
		31: note_dur = CYCLES_PER_US * 781;
		32: note_dur = CYCLES_PER_US * 92969;
		33: note_dur = CYCLES_PER_US * 781;
		34: note_dur = CYCLES_PER_US * 92969;
		35: note_dur = CYCLES_PER_US * 781;
		36: note_dur = CYCLES_PER_US * 374219;
		37: note_dur = CYCLES_PER_US * 781;
		38: note_dur = CYCLES_PER_US * 1124219;
		39: note_dur = CYCLES_PER_US * 781;
		40: note_dur = CYCLES_PER_US * 92969;
		41: note_dur = CYCLES_PER_US * 781;
		42: note_dur = CYCLES_PER_US * 92969;
		43: note_dur = CYCLES_PER_US * 781;
		44: note_dur = CYCLES_PER_US * 92969;
		45: note_dur = CYCLES_PER_US * 781;
		46: note_dur = CYCLES_PER_US * 92969;
		47: note_dur = CYCLES_PER_US * 781;
		48: note_dur = CYCLES_PER_US * 374219;
		49: note_dur = CYCLES_PER_US * 781;
		50: note_dur = CYCLES_PER_US * 1124219;
		51: note_dur = CYCLES_PER_US * 781;
		52: note_dur = CYCLES_PER_US * 186719;
		53: note_dur = CYCLES_PER_US * 781;
		54: note_dur = CYCLES_PER_US * 186719;
		55: note_dur = CYCLES_PER_US * 781;
		56: note_dur = CYCLES_PER_US * 186719;
		57: note_dur = CYCLES_PER_US * 781;
		58: note_dur = CYCLES_PER_US * 186719;
		59: note_dur = CYCLES_PER_US * 781;
		60: note_dur = CYCLES_PER_US * 186719;
		61: note_dur = CYCLES_PER_US * 781;
		62: note_dur = CYCLES_PER_US * 186719;
		63: note_dur = CYCLES_PER_US * 781;
		64: note_dur = CYCLES_PER_US * 186719;
		65: note_dur = CYCLES_PER_US * 781;
		66: note_dur = CYCLES_PER_US * 186719;
		67: note_dur = CYCLES_PER_US * 781;
		68: note_dur = CYCLES_PER_US * 374219;
		69: note_dur = CYCLES_PER_US * 781;
		70: note_dur = CYCLES_PER_US * 186719;
		71: note_dur = CYCLES_PER_US * 781;
		72: note_dur = CYCLES_PER_US * 92969;
		73: note_dur = CYCLES_PER_US * 781;
		74: note_dur = CYCLES_PER_US * 92969;
		75: note_dur = CYCLES_PER_US * 781;
		76: note_dur = CYCLES_PER_US * 374219;
		77: note_dur = CYCLES_PER_US * 781;
		78: note_dur = CYCLES_PER_US * 1124219;
		79: note_dur = CYCLES_PER_US * 781;
		80: note_dur = CYCLES_PER_US * 92969;
		81: note_dur = CYCLES_PER_US * 781;
		82: note_dur = CYCLES_PER_US * 92969;
		83: note_dur = CYCLES_PER_US * 781;
		84: note_dur = CYCLES_PER_US * 92969;
		85: note_dur = CYCLES_PER_US * 781;
		86: note_dur = CYCLES_PER_US * 92969;
		87: note_dur = CYCLES_PER_US * 781;
		88: note_dur = CYCLES_PER_US * 374219;
		89: note_dur = CYCLES_PER_US * 781;
		90: note_dur = CYCLES_PER_US * 1124219;
		91: note_dur = CYCLES_PER_US * 781;
		92: note_dur = CYCLES_PER_US * 92969;
		93: note_dur = CYCLES_PER_US * 781;
		94: note_dur = CYCLES_PER_US * 92969;
		95: note_dur = CYCLES_PER_US * 781;
		96: note_dur = CYCLES_PER_US * 92969;
		97: note_dur = CYCLES_PER_US * 781;
		98: note_dur = CYCLES_PER_US * 92969;
		99: note_dur = CYCLES_PER_US * 781;
		100: note_dur = CYCLES_PER_US * 374219;
		101: note_dur = CYCLES_PER_US * 781;
		102: note_dur = CYCLES_PER_US * 1124219;
		103: note_dur = CYCLES_PER_US * 750781;
		104: note_dur = CYCLES_PER_US * 186719;
		105: note_dur = CYCLES_PER_US * 781;
		106: note_dur = CYCLES_PER_US * 280469;
		107: note_dur = CYCLES_PER_US * 781;
		108: note_dur = CYCLES_PER_US * 186719;
		109: note_dur = CYCLES_PER_US * 781;
		110: note_dur = CYCLES_PER_US * 280469;
		111: note_dur = CYCLES_PER_US * 781;
		112: note_dur = CYCLES_PER_US * 186719;
		113: note_dur = CYCLES_PER_US * 781;
		114: note_dur = CYCLES_PER_US * 186719;
		115: note_dur = CYCLES_PER_US * 781;
		116: note_dur = CYCLES_PER_US * 186719;
		117: note_dur = CYCLES_PER_US * 781;
		118: note_dur = CYCLES_PER_US * 186719;
		119: note_dur = CYCLES_PER_US * 781;
		120: note_dur = CYCLES_PER_US * 186719;
		121: note_dur = CYCLES_PER_US * 781;
		122: note_dur = CYCLES_PER_US * 280469;
		123: note_dur = CYCLES_PER_US * 781;
		124: note_dur = CYCLES_PER_US * 186719;
		125: note_dur = CYCLES_PER_US * 781;
		126: note_dur = CYCLES_PER_US * 280469;
		127: note_dur = CYCLES_PER_US * 781;
		128: note_dur = CYCLES_PER_US * 186719;
		129: note_dur = CYCLES_PER_US * 781;
		130: note_dur = CYCLES_PER_US * 186719;
		131: note_dur = CYCLES_PER_US * 781;
		132: note_dur = CYCLES_PER_US * 186719;
		133: note_dur = CYCLES_PER_US * 781;
		134: note_dur = CYCLES_PER_US * 186719;
		135: note_dur = CYCLES_PER_US * 781;
		136: note_dur = CYCLES_PER_US * 186719;
		137: note_dur = CYCLES_PER_US * 781;
		138: note_dur = CYCLES_PER_US * 280469;
		139: note_dur = CYCLES_PER_US * 781;
		140: note_dur = CYCLES_PER_US * 186719;
		141: note_dur = CYCLES_PER_US * 781;
		142: note_dur = CYCLES_PER_US * 280469;
		143: note_dur = CYCLES_PER_US * 781;
		144: note_dur = CYCLES_PER_US * 186719;
		145: note_dur = CYCLES_PER_US * 781;
		146: note_dur = CYCLES_PER_US * 186719;
		147: note_dur = CYCLES_PER_US * 781;
		148: note_dur = CYCLES_PER_US * 186719;
		149: note_dur = CYCLES_PER_US * 781;
		150: note_dur = CYCLES_PER_US * 186719;
		151: note_dur = CYCLES_PER_US * 781;
		152: note_dur = CYCLES_PER_US * 186719;
		153: note_dur = CYCLES_PER_US * 781;
		154: note_dur = CYCLES_PER_US * 186719;
		155: note_dur = CYCLES_PER_US * 781;
		156: note_dur = CYCLES_PER_US * 186719;
		157: note_dur = CYCLES_PER_US * 781;
		158: note_dur = CYCLES_PER_US * 186719;
		159: note_dur = CYCLES_PER_US * 781;
		160: note_dur = CYCLES_PER_US * 374219;
		161: note_dur = CYCLES_PER_US * 781;
		162: note_dur = CYCLES_PER_US * 186719;
		163: note_dur = CYCLES_PER_US * 781;
		164: note_dur = CYCLES_PER_US * 186719;
		165: note_dur = CYCLES_PER_US * 781;
		166: note_dur = CYCLES_PER_US * 186719;
		167: note_dur = CYCLES_PER_US * 781;
		168: note_dur = CYCLES_PER_US * 186719;
		169: note_dur = CYCLES_PER_US * 781;
		170: note_dur = CYCLES_PER_US * 186719;
		171: note_dur = CYCLES_PER_US * 781;
		172: note_dur = CYCLES_PER_US * 280469;
		173: note_dur = CYCLES_PER_US * 781;
		174: note_dur = CYCLES_PER_US * 186719;
		175: note_dur = CYCLES_PER_US * 781;
		176: note_dur = CYCLES_PER_US * 280469;
		177: note_dur = CYCLES_PER_US * 781;
		178: note_dur = CYCLES_PER_US * 186719;
		179: note_dur = CYCLES_PER_US * 781;
		180: note_dur = CYCLES_PER_US * 280469;
		181: note_dur = CYCLES_PER_US * 781;
		182: note_dur = CYCLES_PER_US * 186719;
		183: note_dur = CYCLES_PER_US * 781;
		184: note_dur = CYCLES_PER_US * 186719;
		185: note_dur = CYCLES_PER_US * 781;
		186: note_dur = CYCLES_PER_US * 280469;
		187: note_dur = CYCLES_PER_US * 781;
		188: note_dur = CYCLES_PER_US * 186719;
		189: note_dur = CYCLES_PER_US * 781;
		190: note_dur = CYCLES_PER_US * 280469;
		191: note_dur = CYCLES_PER_US * 781;
		192: note_dur = CYCLES_PER_US * 186719;
		193: note_dur = CYCLES_PER_US * 781;
		194: note_dur = CYCLES_PER_US * 186719;
		195: note_dur = CYCLES_PER_US * 781;
		196: note_dur = CYCLES_PER_US * 186719;
		197: note_dur = CYCLES_PER_US * 781;
		198: note_dur = CYCLES_PER_US * 186719;
		199: note_dur = CYCLES_PER_US * 781;
		200: note_dur = CYCLES_PER_US * 186719;
		201: note_dur = CYCLES_PER_US * 781;
		202: note_dur = CYCLES_PER_US * 280469;
		203: note_dur = CYCLES_PER_US * 781;
		204: note_dur = CYCLES_PER_US * 186719;
		205: note_dur = CYCLES_PER_US * 781;
		206: note_dur = CYCLES_PER_US * 280469;
		207: note_dur = CYCLES_PER_US * 781;
		208: note_dur = CYCLES_PER_US * 186719;
		209: note_dur = CYCLES_PER_US * 781;
		210: note_dur = CYCLES_PER_US * 186719;
		211: note_dur = CYCLES_PER_US * 781;
		212: note_dur = CYCLES_PER_US * 186719;
		213: note_dur = CYCLES_PER_US * 781;
		214: note_dur = CYCLES_PER_US * 186719;
		215: note_dur = CYCLES_PER_US * 781;
		216: note_dur = CYCLES_PER_US * 1124219;
		217: note_dur = CYCLES_PER_US * 0;
		218: note_dur = CYCLES_PER_US * 186719;
		219: note_dur = CYCLES_PER_US * 781;
		220: note_dur = CYCLES_PER_US * 186719;
		221: note_dur = CYCLES_PER_US * 781;
		222: note_dur = CYCLES_PER_US * 186719;
		223: note_dur = CYCLES_PER_US * 781;
		224: note_dur = CYCLES_PER_US * 186719;
		225: note_dur = CYCLES_PER_US * 781;
		226: note_dur = CYCLES_PER_US * 186719;
		227: note_dur = CYCLES_PER_US * 781;
		228: note_dur = CYCLES_PER_US * 186719;
		229: note_dur = CYCLES_PER_US * 781;
		230: note_dur = CYCLES_PER_US * 186719;
		231: note_dur = CYCLES_PER_US * 781;
		232: note_dur = CYCLES_PER_US * 186719;
		233: note_dur = CYCLES_PER_US * 781;
		234: note_dur = CYCLES_PER_US * 374219;
		235: note_dur = CYCLES_PER_US * 781;
		236: note_dur = CYCLES_PER_US * 186719;
		237: note_dur = CYCLES_PER_US * 781;
		238: note_dur = CYCLES_PER_US * 92969;
		239: note_dur = CYCLES_PER_US * 781;
		240: note_dur = CYCLES_PER_US * 92969;
		241: note_dur = CYCLES_PER_US * 781;
		242: note_dur = CYCLES_PER_US * 374219;
		243: note_dur = CYCLES_PER_US * 781;
		244: note_dur = CYCLES_PER_US * 1124219;
		245: note_dur = CYCLES_PER_US * 781;
		246: note_dur = CYCLES_PER_US * 92969;
		247: note_dur = CYCLES_PER_US * 781;
		248: note_dur = CYCLES_PER_US * 92969;
		249: note_dur = CYCLES_PER_US * 781;
		250: note_dur = CYCLES_PER_US * 92969;
		251: note_dur = CYCLES_PER_US * 781;
		252: note_dur = CYCLES_PER_US * 92969;
		253: note_dur = CYCLES_PER_US * 781;
		254: note_dur = CYCLES_PER_US * 374219;
		255: note_dur = CYCLES_PER_US * 781;
		256: note_dur = CYCLES_PER_US * 1124219;
		257: note_dur = CYCLES_PER_US * 781;
		258: note_dur = CYCLES_PER_US * 92969;
		259: note_dur = CYCLES_PER_US * 781;
		260: note_dur = CYCLES_PER_US * 92969;
		261: note_dur = CYCLES_PER_US * 781;
		262: note_dur = CYCLES_PER_US * 92969;
		263: note_dur = CYCLES_PER_US * 781;
		264: note_dur = CYCLES_PER_US * 92969;
		265: note_dur = CYCLES_PER_US * 781;
		266: note_dur = CYCLES_PER_US * 374219;
		267: note_dur = CYCLES_PER_US * 781;
		268: note_dur = CYCLES_PER_US * 1124219;
		269: note_dur = CYCLES_PER_US * 781;
		270: note_dur = CYCLES_PER_US * 186719;
		271: note_dur = CYCLES_PER_US * 781;
		272: note_dur = CYCLES_PER_US * 186719;
		273: note_dur = CYCLES_PER_US * 781;
		274: note_dur = CYCLES_PER_US * 186719;
		275: note_dur = CYCLES_PER_US * 781;
		276: note_dur = CYCLES_PER_US * 186719;
		277: note_dur = CYCLES_PER_US * 781;
		278: note_dur = CYCLES_PER_US * 186719;
		279: note_dur = CYCLES_PER_US * 781;
		280: note_dur = CYCLES_PER_US * 186719;
		281: note_dur = CYCLES_PER_US * 781;
		282: note_dur = CYCLES_PER_US * 186719;
		283: note_dur = CYCLES_PER_US * 781;
		284: note_dur = CYCLES_PER_US * 186719;
		285: note_dur = CYCLES_PER_US * 781;
		286: note_dur = CYCLES_PER_US * 374219;
		287: note_dur = CYCLES_PER_US * 781;
		288: note_dur = CYCLES_PER_US * 186719;
		289: note_dur = CYCLES_PER_US * 781;
		290: note_dur = CYCLES_PER_US * 92969;
		291: note_dur = CYCLES_PER_US * 781;
		292: note_dur = CYCLES_PER_US * 92969;
		293: note_dur = CYCLES_PER_US * 781;
		294: note_dur = CYCLES_PER_US * 374219;
		295: note_dur = CYCLES_PER_US * 781;
		296: note_dur = CYCLES_PER_US * 1124219;
		297: note_dur = CYCLES_PER_US * 781;
		298: note_dur = CYCLES_PER_US * 92969;
		299: note_dur = CYCLES_PER_US * 781;
		300: note_dur = CYCLES_PER_US * 92969;
		301: note_dur = CYCLES_PER_US * 781;
		302: note_dur = CYCLES_PER_US * 92969;
		303: note_dur = CYCLES_PER_US * 781;
		304: note_dur = CYCLES_PER_US * 92969;
		305: note_dur = CYCLES_PER_US * 781;
		306: note_dur = CYCLES_PER_US * 374219;
		307: note_dur = CYCLES_PER_US * 781;
		308: note_dur = CYCLES_PER_US * 1124219;
		309: note_dur = CYCLES_PER_US * 781;
		310: note_dur = CYCLES_PER_US * 92969;
		311: note_dur = CYCLES_PER_US * 781;
		312: note_dur = CYCLES_PER_US * 92969;
		313: note_dur = CYCLES_PER_US * 781;
		314: note_dur = CYCLES_PER_US * 92969;
		315: note_dur = CYCLES_PER_US * 781;
		316: note_dur = CYCLES_PER_US * 92969;
		317: note_dur = CYCLES_PER_US * 781;
		318: note_dur = CYCLES_PER_US * 374219;
		319: note_dur = CYCLES_PER_US * 781;
		320: note_dur = CYCLES_PER_US * 1124219;
		321: note_dur = CYCLES_PER_US * 563281;
		322: note_dur = CYCLES_PER_US * 0;
		323: note_dur = CYCLES_PER_US * 749219;
		324: note_dur = CYCLES_PER_US * 187500;
		325: note_dur = CYCLES_PER_US * 781;
		326: note_dur = CYCLES_PER_US * 92969;
		327: note_dur = CYCLES_PER_US * 781;
		328: note_dur = CYCLES_PER_US * 92969;
		329: note_dur = CYCLES_PER_US * 781;
		330: note_dur = CYCLES_PER_US * 749219;
		331: note_dur = CYCLES_PER_US * 781;
		332: note_dur = CYCLES_PER_US * 561719;
		333: note_dur = CYCLES_PER_US * 781;
		334: note_dur = CYCLES_PER_US * 186719;
		335: note_dur = CYCLES_PER_US * 781;
		336: note_dur = CYCLES_PER_US * 374219;
		337: note_dur = CYCLES_PER_US * 750781;
		338: note_dur = CYCLES_PER_US * 186719;
		339: note_dur = CYCLES_PER_US * 781;
		340: note_dur = CYCLES_PER_US * 186719;
		341: note_dur = CYCLES_PER_US * 781;
		342: note_dur = CYCLES_PER_US * 186719;
		343: note_dur = CYCLES_PER_US * 781;
		344: note_dur = CYCLES_PER_US * 186719;
		345: note_dur = CYCLES_PER_US * 781;
		346: note_dur = CYCLES_PER_US * 186719;
		347: note_dur = CYCLES_PER_US * 781;
		348: note_dur = CYCLES_PER_US * 561719;
		349: note_dur = CYCLES_PER_US * 781;
		350: note_dur = CYCLES_PER_US * 374219;
		351: note_dur = CYCLES_PER_US * 781;
		352: note_dur = CYCLES_PER_US * 561719;
		353: note_dur = CYCLES_PER_US * 781;
		354: note_dur = CYCLES_PER_US * 186719;
		355: note_dur = CYCLES_PER_US * 781;
		356: note_dur = CYCLES_PER_US * 186719;
		357: note_dur = CYCLES_PER_US * 781;
		358: note_dur = CYCLES_PER_US * 92969;
		359: note_dur = CYCLES_PER_US * 750781;
		360: note_dur = CYCLES_PER_US * 561719;
		361: note_dur = CYCLES_PER_US * 781;
		362: note_dur = CYCLES_PER_US * 280469;
		363: note_dur = CYCLES_PER_US * 781;
		364: note_dur = CYCLES_PER_US * 186719;
		365: note_dur = CYCLES_PER_US * 781;
		366: note_dur = CYCLES_PER_US * 374219;
		367: note_dur = CYCLES_PER_US * 781;
		368: note_dur = CYCLES_PER_US * 280469;
		369: note_dur = CYCLES_PER_US * 781;
		370: note_dur = CYCLES_PER_US * 561719;
		371: note_dur = CYCLES_PER_US * 781;
		372: note_dur = CYCLES_PER_US * 280469;
		373: note_dur = CYCLES_PER_US * 781;
		374: note_dur = CYCLES_PER_US * 186719;
		375: note_dur = CYCLES_PER_US * 781;
		376: note_dur = CYCLES_PER_US * 186719;
		377: note_dur = CYCLES_PER_US * 781;
		378: note_dur = CYCLES_PER_US * 186719;
		379: note_dur = CYCLES_PER_US * 781;
		380: note_dur = CYCLES_PER_US * 186719;
		381: note_dur = CYCLES_PER_US * 781;
		382: note_dur = CYCLES_PER_US * 186719;
		383: note_dur = CYCLES_PER_US * 781;
		384: note_dur = CYCLES_PER_US * 561719;
		385: note_dur = CYCLES_PER_US * 781;
		386: note_dur = CYCLES_PER_US * 280469;
		387: note_dur = CYCLES_PER_US * 781;
		388: note_dur = CYCLES_PER_US * 186719;
		389: note_dur = CYCLES_PER_US * 781;
		390: note_dur = CYCLES_PER_US * 374219;
		391: note_dur = CYCLES_PER_US * 781;
		392: note_dur = CYCLES_PER_US * 280469;
		393: note_dur = CYCLES_PER_US * 781;
		394: note_dur = CYCLES_PER_US * 561719;
		395: note_dur = CYCLES_PER_US * 781;
		396: note_dur = CYCLES_PER_US * 280469;
		397: note_dur = CYCLES_PER_US * 781;
		398: note_dur = CYCLES_PER_US * 186719;
		399: note_dur = CYCLES_PER_US * 781;
		400: note_dur = CYCLES_PER_US * 186719;
		401: note_dur = CYCLES_PER_US * 781;
		402: note_dur = CYCLES_PER_US * 92969;
		403: note_dur = CYCLES_PER_US * 563281;
		404: note_dur = CYCLES_PER_US * 1311719;
		405: note_dur = CYCLES_PER_US * 563281;
		406: note_dur = CYCLES_PER_US * 186719;
		407: note_dur = CYCLES_PER_US * 188281;
		408: note_dur = CYCLES_PER_US * 186719;
		409: note_dur = CYCLES_PER_US * 781;
		410: note_dur = CYCLES_PER_US * 749219;
		411: note_dur = CYCLES_PER_US * 781;
		412: note_dur = CYCLES_PER_US * 374219;
		413: note_dur = CYCLES_PER_US * 781;
		414: note_dur = CYCLES_PER_US * 1124219;
		415: note_dur = CYCLES_PER_US * 188281;
		416: note_dur = CYCLES_PER_US * 186719;
		417: note_dur = CYCLES_PER_US * 781;
		418: note_dur = CYCLES_PER_US * 186719;
		419: note_dur = CYCLES_PER_US * 781;
		420: note_dur = CYCLES_PER_US * 186719;
		421: note_dur = CYCLES_PER_US * 188281;
		422: note_dur = CYCLES_PER_US * 936719;
		423: note_dur = CYCLES_PER_US * 375781;
		424: note_dur = CYCLES_PER_US * 374219;
		425: note_dur = CYCLES_PER_US * 781;
		426: note_dur = CYCLES_PER_US * 561719;
		427: note_dur = CYCLES_PER_US * 781;
		428: note_dur = CYCLES_PER_US * 186719;
		429: note_dur = CYCLES_PER_US * 375781;
		430: note_dur = CYCLES_PER_US * 374219;
		431: note_dur = CYCLES_PER_US * 781;
		432: note_dur = CYCLES_PER_US * 374219;
		433: note_dur = CYCLES_PER_US * 781;
		434: note_dur = CYCLES_PER_US * 561719;
		435: note_dur = CYCLES_PER_US * 781;
		436: note_dur = CYCLES_PER_US * 374219;
		437: note_dur = CYCLES_PER_US * 781;
		438: note_dur = CYCLES_PER_US * 186719;
		439: note_dur = CYCLES_PER_US * 781;
		440: note_dur = CYCLES_PER_US * 186719;
		441: note_dur = CYCLES_PER_US * 781;
		442: note_dur = CYCLES_PER_US * 186719;
		443: note_dur = CYCLES_PER_US * 781;
		444: note_dur = CYCLES_PER_US * 186719;
		445: note_dur = CYCLES_PER_US * 781;
		446: note_dur = CYCLES_PER_US * 186719;
		447: note_dur = CYCLES_PER_US * 781;
		448: note_dur = CYCLES_PER_US * 561719;
		449: note_dur = CYCLES_PER_US * 781;
		450: note_dur = CYCLES_PER_US * 374219;
		451: note_dur = CYCLES_PER_US * 781;
		452: note_dur = CYCLES_PER_US * 186719;
		453: note_dur = CYCLES_PER_US * 781;
		454: note_dur = CYCLES_PER_US * 374219;
		455: note_dur = CYCLES_PER_US * 781;
		456: note_dur = CYCLES_PER_US * 280469;
		457: note_dur = CYCLES_PER_US * 781;
		458: note_dur = CYCLES_PER_US * 561719;
		459: note_dur = CYCLES_PER_US * 781;
		460: note_dur = CYCLES_PER_US * 374219;
		461: note_dur = CYCLES_PER_US * 781;
		462: note_dur = CYCLES_PER_US * 186719;
		463: note_dur = CYCLES_PER_US * 781;
		464: note_dur = CYCLES_PER_US * 186719;
		465: note_dur = CYCLES_PER_US * 781;
		466: note_dur = CYCLES_PER_US * 186719;
		467: note_dur = CYCLES_PER_US * 781;
		468: note_dur = CYCLES_PER_US * 186719;
		469: note_dur = CYCLES_PER_US * 781;
		470: note_dur = CYCLES_PER_US * 0;
		471: note_dur = CYCLES_PER_US * 186719;
		472: note_dur = CYCLES_PER_US * 0;
		473: note_dur = CYCLES_PER_US * 93750;
		474: note_dur = CYCLES_PER_US * 0;
		475: note_dur = CYCLES_PER_US * 92969;
		476: note_dur = CYCLES_PER_US * 0;
		477: note_dur = CYCLES_PER_US * 186719;
		478: note_dur = CYCLES_PER_US * 562500;
		479: note_dur = CYCLES_PER_US * 781;
		480: note_dur = CYCLES_PER_US * 92969;
		481: note_dur = CYCLES_PER_US * 781;
		482: note_dur = CYCLES_PER_US * 92969;
		483: note_dur = CYCLES_PER_US * 781;
		484: note_dur = CYCLES_PER_US * 374219;
		485: note_dur = CYCLES_PER_US * 375781;
		486: note_dur = CYCLES_PER_US * 561719;
		487: note_dur = CYCLES_PER_US * 781;
		488: note_dur = CYCLES_PER_US * 186719;
		489: note_dur = CYCLES_PER_US * 781;
		490: note_dur = CYCLES_PER_US * 374219;
		491: note_dur = CYCLES_PER_US * 750781;
		492: note_dur = CYCLES_PER_US * 561719;
		493: note_dur = CYCLES_PER_US * 781;
		494: note_dur = CYCLES_PER_US * 92969;
		495: note_dur = CYCLES_PER_US * 781;
		496: note_dur = CYCLES_PER_US * 92969;
		497: note_dur = CYCLES_PER_US * 781;
		498: note_dur = CYCLES_PER_US * 186719;
		499: note_dur = CYCLES_PER_US * 781;
		500: note_dur = CYCLES_PER_US * 186719;
		501: note_dur = CYCLES_PER_US * 781;
		502: note_dur = CYCLES_PER_US * 186719;
		503: note_dur = CYCLES_PER_US * 781;
		504: note_dur = CYCLES_PER_US * 186719;
		505: note_dur = CYCLES_PER_US * 781;
		506: note_dur = CYCLES_PER_US * 186719;
		507: note_dur = CYCLES_PER_US * 781;
		508: note_dur = CYCLES_PER_US * 186719;
		509: note_dur = CYCLES_PER_US * 781;
		510: note_dur = CYCLES_PER_US * 186719;
		511: note_dur = CYCLES_PER_US * 781;
		512: note_dur = CYCLES_PER_US * 561719;
		513: note_dur = CYCLES_PER_US * 781;
		514: note_dur = CYCLES_PER_US * 374219;
		515: note_dur = CYCLES_PER_US * 750781;
		516: note_dur = CYCLES_PER_US * 561719;
		517: note_dur = CYCLES_PER_US * 781;
		518: note_dur = CYCLES_PER_US * 186719;
		519: note_dur = CYCLES_PER_US * 188281;
		520: note_dur = CYCLES_PER_US * 186719;
		521: note_dur = CYCLES_PER_US * 781;
		522: note_dur = CYCLES_PER_US * 186719;
		523: note_dur = CYCLES_PER_US * 781;
		524: note_dur = CYCLES_PER_US * 186719;
		525: note_dur = CYCLES_PER_US * 781;
		526: note_dur = CYCLES_PER_US * 374219;
		527: note_dur = CYCLES_PER_US * 781;
		528: note_dur = CYCLES_PER_US * 561719;
		529: note_dur = CYCLES_PER_US * 781;
		530: note_dur = CYCLES_PER_US * 186719;
		531: note_dur = CYCLES_PER_US * 375781;
		532: note_dur = CYCLES_PER_US * 186719;
		533: note_dur = CYCLES_PER_US * 781;
		534: note_dur = CYCLES_PER_US * 186719;
		535: note_dur = CYCLES_PER_US * 781;
		536: note_dur = CYCLES_PER_US * 374219;
		537: note_dur = CYCLES_PER_US * 781;
		538: note_dur = CYCLES_PER_US * 561719;
		539: note_dur = CYCLES_PER_US * 781;
		540: note_dur = CYCLES_PER_US * 186719;
		541: note_dur = CYCLES_PER_US * 188281;
		542: note_dur = CYCLES_PER_US * 186719;
		543: note_dur = CYCLES_PER_US * 781;
		544: note_dur = CYCLES_PER_US * 186719;
		545: note_dur = CYCLES_PER_US * 781;
		546: note_dur = CYCLES_PER_US * 186719;
		547: note_dur = CYCLES_PER_US * 781;
		548: note_dur = CYCLES_PER_US * 374219;
		549: note_dur = CYCLES_PER_US * 781;
		550: note_dur = CYCLES_PER_US * 561719;
		551: note_dur = CYCLES_PER_US * 781;
		552: note_dur = CYCLES_PER_US * 374219;
		553: note_dur = CYCLES_PER_US * 781;
		554: note_dur = CYCLES_PER_US * 186719;
		555: note_dur = CYCLES_PER_US * 781;
		556: note_dur = CYCLES_PER_US * 561719;
		557: note_dur = CYCLES_PER_US * 781;
		558: note_dur = CYCLES_PER_US * 186719;
		559: note_dur = CYCLES_PER_US * 781;
		560: note_dur = CYCLES_PER_US * 2249219;
		561: note_dur = CYCLES_PER_US * 19500781;
		562: note_dur = CYCLES_PER_US * 186719;
		563: note_dur = CYCLES_PER_US * 781;
		564: note_dur = CYCLES_PER_US * 186719;
		565: note_dur = CYCLES_PER_US * 781;
		566: note_dur = CYCLES_PER_US * 186719;
		567: note_dur = CYCLES_PER_US * 781;
		568: note_dur = CYCLES_PER_US * 186719;
		569: note_dur = CYCLES_PER_US * 781;
		570: note_dur = CYCLES_PER_US * 2249219;
		571: note_dur = CYCLES_PER_US * 19500781;
		572: note_dur = CYCLES_PER_US * 186719;
		573: note_dur = CYCLES_PER_US * 781;
		574: note_dur = CYCLES_PER_US * 186719;
		575: note_dur = CYCLES_PER_US * 781;
		576: note_dur = CYCLES_PER_US * 186719;
		577: note_dur = CYCLES_PER_US * 781;
		578: note_dur = CYCLES_PER_US * 186719;
		579: note_dur = CYCLES_PER_US * 781;
		580: note_dur = CYCLES_PER_US * 186719;
		581: note_dur = CYCLES_PER_US * 781;
		582: note_dur = CYCLES_PER_US * 186719;
		583: note_dur = CYCLES_PER_US * 781;
		584: note_dur = CYCLES_PER_US * 186719;
		585: note_dur = CYCLES_PER_US * 781;
		586: note_dur = CYCLES_PER_US * 186719;
		587: note_dur = CYCLES_PER_US * 781;
		588: note_dur = CYCLES_PER_US * 374219;
		589: note_dur = CYCLES_PER_US * 781;
		590: note_dur = CYCLES_PER_US * 186719;
		591: note_dur = CYCLES_PER_US * 781;
		592: note_dur = CYCLES_PER_US * 92969;
		593: note_dur = CYCLES_PER_US * 781;
		594: note_dur = CYCLES_PER_US * 92969;
		595: note_dur = CYCLES_PER_US * 781;
		596: note_dur = CYCLES_PER_US * 374219;
		597: note_dur = CYCLES_PER_US * 781;
		598: note_dur = CYCLES_PER_US * 1124219;
		599: note_dur = CYCLES_PER_US * 781;
		600: note_dur = CYCLES_PER_US * 92969;
		601: note_dur = CYCLES_PER_US * 781;
		602: note_dur = CYCLES_PER_US * 92969;
		603: note_dur = CYCLES_PER_US * 781;
		604: note_dur = CYCLES_PER_US * 92969;
		605: note_dur = CYCLES_PER_US * 781;
		606: note_dur = CYCLES_PER_US * 92969;
		607: note_dur = CYCLES_PER_US * 781;
		608: note_dur = CYCLES_PER_US * 374219;
		609: note_dur = CYCLES_PER_US * 781;
		610: note_dur = CYCLES_PER_US * 1124219;
		611: note_dur = CYCLES_PER_US * 781;
		612: note_dur = CYCLES_PER_US * 92969;
		613: note_dur = CYCLES_PER_US * 781;
		614: note_dur = CYCLES_PER_US * 92969;
		615: note_dur = CYCLES_PER_US * 781;
		616: note_dur = CYCLES_PER_US * 92969;
		617: note_dur = CYCLES_PER_US * 781;
		618: note_dur = CYCLES_PER_US * 92969;
		619: note_dur = CYCLES_PER_US * 781;
		620: note_dur = CYCLES_PER_US * 374219;
		621: note_dur = CYCLES_PER_US * 781;
		622: note_dur = CYCLES_PER_US * 1124219;
		623: note_dur = CYCLES_PER_US * 781;
		624: note_dur = CYCLES_PER_US * 186719;
		625: note_dur = CYCLES_PER_US * 781;
		626: note_dur = CYCLES_PER_US * 186719;
		627: note_dur = CYCLES_PER_US * 781;
		628: note_dur = CYCLES_PER_US * 186719;
		629: note_dur = CYCLES_PER_US * 781;
		630: note_dur = CYCLES_PER_US * 186719;
		631: note_dur = CYCLES_PER_US * 781;
		632: note_dur = CYCLES_PER_US * 186719;
		633: note_dur = CYCLES_PER_US * 781;
		634: note_dur = CYCLES_PER_US * 186719;
		635: note_dur = CYCLES_PER_US * 781;
		636: note_dur = CYCLES_PER_US * 186719;
		637: note_dur = CYCLES_PER_US * 781;
		638: note_dur = CYCLES_PER_US * 186719;
		639: note_dur = CYCLES_PER_US * 781;
		640: note_dur = CYCLES_PER_US * 374219;
		641: note_dur = CYCLES_PER_US * 781;
		642: note_dur = CYCLES_PER_US * 186719;
		643: note_dur = CYCLES_PER_US * 781;
		644: note_dur = CYCLES_PER_US * 92969;
		645: note_dur = CYCLES_PER_US * 781;
		646: note_dur = CYCLES_PER_US * 92969;
		647: note_dur = CYCLES_PER_US * 781;
		648: note_dur = CYCLES_PER_US * 374219;
		649: note_dur = CYCLES_PER_US * 781;
		650: note_dur = CYCLES_PER_US * 1124219;
		651: note_dur = CYCLES_PER_US * 781;
		652: note_dur = CYCLES_PER_US * 92969;
		653: note_dur = CYCLES_PER_US * 781;
		654: note_dur = CYCLES_PER_US * 92969;
		655: note_dur = CYCLES_PER_US * 781;
		656: note_dur = CYCLES_PER_US * 92969;
		657: note_dur = CYCLES_PER_US * 781;
		658: note_dur = CYCLES_PER_US * 92969;
		659: note_dur = CYCLES_PER_US * 781;
		660: note_dur = CYCLES_PER_US * 374219;
		661: note_dur = CYCLES_PER_US * 781;
		662: note_dur = CYCLES_PER_US * 1124219;
		663: note_dur = CYCLES_PER_US * 781;
		664: note_dur = CYCLES_PER_US * 92969;
		665: note_dur = CYCLES_PER_US * 781;
		666: note_dur = CYCLES_PER_US * 92969;
		667: note_dur = CYCLES_PER_US * 781;
		668: note_dur = CYCLES_PER_US * 92969;
		669: note_dur = CYCLES_PER_US * 781;
		670: note_dur = CYCLES_PER_US * 92969;
		671: note_dur = CYCLES_PER_US * 781;
		672: note_dur = CYCLES_PER_US * 374219;
		673: note_dur = CYCLES_PER_US * 781;
		674: note_dur = CYCLES_PER_US * 1124219;
		675: note_dur = CYCLES_PER_US * 750781;
		676: note_dur = CYCLES_PER_US * 186719;
		677: note_dur = CYCLES_PER_US * 781;
		678: note_dur = CYCLES_PER_US * 280469;
		679: note_dur = CYCLES_PER_US * 781;
		680: note_dur = CYCLES_PER_US * 186719;
		681: note_dur = CYCLES_PER_US * 781;
		682: note_dur = CYCLES_PER_US * 280469;
		683: note_dur = CYCLES_PER_US * 781;
		684: note_dur = CYCLES_PER_US * 186719;
		685: note_dur = CYCLES_PER_US * 781;
		686: note_dur = CYCLES_PER_US * 186719;
		687: note_dur = CYCLES_PER_US * 781;
		688: note_dur = CYCLES_PER_US * 186719;
		689: note_dur = CYCLES_PER_US * 781;
		690: note_dur = CYCLES_PER_US * 186719;
		691: note_dur = CYCLES_PER_US * 781;
		692: note_dur = CYCLES_PER_US * 186719;
		693: note_dur = CYCLES_PER_US * 781;
		694: note_dur = CYCLES_PER_US * 280469;
		695: note_dur = CYCLES_PER_US * 781;
		696: note_dur = CYCLES_PER_US * 186719;
		697: note_dur = CYCLES_PER_US * 781;
		698: note_dur = CYCLES_PER_US * 280469;
		699: note_dur = CYCLES_PER_US * 781;
		700: note_dur = CYCLES_PER_US * 186719;
		701: note_dur = CYCLES_PER_US * 781;
		702: note_dur = CYCLES_PER_US * 186719;
		703: note_dur = CYCLES_PER_US * 781;
		704: note_dur = CYCLES_PER_US * 186719;
		705: note_dur = CYCLES_PER_US * 781;
		706: note_dur = CYCLES_PER_US * 186719;
		707: note_dur = CYCLES_PER_US * 781;
		708: note_dur = CYCLES_PER_US * 186719;
		709: note_dur = CYCLES_PER_US * 781;
		710: note_dur = CYCLES_PER_US * 280469;
		711: note_dur = CYCLES_PER_US * 781;
		712: note_dur = CYCLES_PER_US * 186719;
		713: note_dur = CYCLES_PER_US * 781;
		714: note_dur = CYCLES_PER_US * 280469;
		715: note_dur = CYCLES_PER_US * 781;
		716: note_dur = CYCLES_PER_US * 186719;
		717: note_dur = CYCLES_PER_US * 781;
		718: note_dur = CYCLES_PER_US * 186719;
		719: note_dur = CYCLES_PER_US * 781;
		720: note_dur = CYCLES_PER_US * 186719;
		721: note_dur = CYCLES_PER_US * 781;
		722: note_dur = CYCLES_PER_US * 186719;
		723: note_dur = CYCLES_PER_US * 781;
		724: note_dur = CYCLES_PER_US * 186719;
		725: note_dur = CYCLES_PER_US * 781;
		726: note_dur = CYCLES_PER_US * 186719;
		727: note_dur = CYCLES_PER_US * 781;
		728: note_dur = CYCLES_PER_US * 186719;
		729: note_dur = CYCLES_PER_US * 781;
		730: note_dur = CYCLES_PER_US * 186719;
		731: note_dur = CYCLES_PER_US * 781;
		732: note_dur = CYCLES_PER_US * 374219;
		733: note_dur = CYCLES_PER_US * 781;
		734: note_dur = CYCLES_PER_US * 186719;
		735: note_dur = CYCLES_PER_US * 781;
		736: note_dur = CYCLES_PER_US * 186719;
		737: note_dur = CYCLES_PER_US * 781;
		738: note_dur = CYCLES_PER_US * 186719;
		739: note_dur = CYCLES_PER_US * 781;
		740: note_dur = CYCLES_PER_US * 186719;
		741: note_dur = CYCLES_PER_US * 781;
		742: note_dur = CYCLES_PER_US * 186719;
		743: note_dur = CYCLES_PER_US * 781;
		744: note_dur = CYCLES_PER_US * 280469;
		745: note_dur = CYCLES_PER_US * 781;
		746: note_dur = CYCLES_PER_US * 186719;
		747: note_dur = CYCLES_PER_US * 781;
		748: note_dur = CYCLES_PER_US * 280469;
		749: note_dur = CYCLES_PER_US * 781;
		750: note_dur = CYCLES_PER_US * 186719;
		751: note_dur = CYCLES_PER_US * 781;
		752: note_dur = CYCLES_PER_US * 280469;
		753: note_dur = CYCLES_PER_US * 781;
		754: note_dur = CYCLES_PER_US * 186719;
		755: note_dur = CYCLES_PER_US * 781;
		756: note_dur = CYCLES_PER_US * 186719;
		757: note_dur = CYCLES_PER_US * 781;
		758: note_dur = CYCLES_PER_US * 280469;
		759: note_dur = CYCLES_PER_US * 781;
		760: note_dur = CYCLES_PER_US * 186719;
		761: note_dur = CYCLES_PER_US * 781;
		762: note_dur = CYCLES_PER_US * 280469;
		763: note_dur = CYCLES_PER_US * 781;
		764: note_dur = CYCLES_PER_US * 186719;
		765: note_dur = CYCLES_PER_US * 781;
		766: note_dur = CYCLES_PER_US * 186719;
		767: note_dur = CYCLES_PER_US * 781;
		768: note_dur = CYCLES_PER_US * 186719;
		769: note_dur = CYCLES_PER_US * 781;
		770: note_dur = CYCLES_PER_US * 186719;
		771: note_dur = CYCLES_PER_US * 781;
		772: note_dur = CYCLES_PER_US * 186719;
		773: note_dur = CYCLES_PER_US * 781;
		774: note_dur = CYCLES_PER_US * 280469;
		775: note_dur = CYCLES_PER_US * 781;
		776: note_dur = CYCLES_PER_US * 186719;
		777: note_dur = CYCLES_PER_US * 781;
		778: note_dur = CYCLES_PER_US * 280469;
		779: note_dur = CYCLES_PER_US * 781;
		780: note_dur = CYCLES_PER_US * 186719;
		781: note_dur = CYCLES_PER_US * 781;
		782: note_dur = CYCLES_PER_US * 186719;
		783: note_dur = CYCLES_PER_US * 781;
		784: note_dur = CYCLES_PER_US * 186719;
		785: note_dur = CYCLES_PER_US * 781;
		786: note_dur = CYCLES_PER_US * 186719;
		787: note_dur = CYCLES_PER_US * 781;
		788: note_dur = CYCLES_PER_US * 1124219;
		789: note_dur = CYCLES_PER_US * 781;
		790: note_dur = CYCLES_PER_US * 186719;
		791: note_dur = CYCLES_PER_US * 781;
		792: note_dur = CYCLES_PER_US * 186719;
		793: note_dur = CYCLES_PER_US * 781;
		794: note_dur = CYCLES_PER_US * 186719;
		795: note_dur = CYCLES_PER_US * 781;
		796: note_dur = CYCLES_PER_US * 186719;
		797: note_dur = CYCLES_PER_US * 781;
		798: note_dur = CYCLES_PER_US * 186719;
		799: note_dur = CYCLES_PER_US * 781;
		800: note_dur = CYCLES_PER_US * 186719;
		801: note_dur = CYCLES_PER_US * 781;
		802: note_dur = CYCLES_PER_US * 186719;
		803: note_dur = CYCLES_PER_US * 781;
		804: note_dur = CYCLES_PER_US * 186719;
		805: note_dur = CYCLES_PER_US * 781;
		806: note_dur = CYCLES_PER_US * 374219;
		807: note_dur = CYCLES_PER_US * 781;
		808: note_dur = CYCLES_PER_US * 186719;
		809: note_dur = CYCLES_PER_US * 781;
		810: note_dur = CYCLES_PER_US * 92969;
		811: note_dur = CYCLES_PER_US * 781;
		812: note_dur = CYCLES_PER_US * 92969;
		813: note_dur = CYCLES_PER_US * 781;
		814: note_dur = CYCLES_PER_US * 374219;
		815: note_dur = CYCLES_PER_US * 781;
		816: note_dur = CYCLES_PER_US * 1124219;
		817: note_dur = CYCLES_PER_US * 781;
		818: note_dur = CYCLES_PER_US * 92969;
		819: note_dur = CYCLES_PER_US * 781;
		820: note_dur = CYCLES_PER_US * 92969;
		821: note_dur = CYCLES_PER_US * 781;
		822: note_dur = CYCLES_PER_US * 92969;
		823: note_dur = CYCLES_PER_US * 781;
		824: note_dur = CYCLES_PER_US * 92969;
		825: note_dur = CYCLES_PER_US * 781;
		826: note_dur = CYCLES_PER_US * 374219;
		827: note_dur = CYCLES_PER_US * 781;
		828: note_dur = CYCLES_PER_US * 1124219;
		829: note_dur = CYCLES_PER_US * 781;
		830: note_dur = CYCLES_PER_US * 92969;
		831: note_dur = CYCLES_PER_US * 781;
		832: note_dur = CYCLES_PER_US * 92969;
		833: note_dur = CYCLES_PER_US * 781;
		834: note_dur = CYCLES_PER_US * 92969;
		835: note_dur = CYCLES_PER_US * 781;
		836: note_dur = CYCLES_PER_US * 92969;
		837: note_dur = CYCLES_PER_US * 781;
		838: note_dur = CYCLES_PER_US * 374219;
		839: note_dur = CYCLES_PER_US * 781;
		840: note_dur = CYCLES_PER_US * 1124219;
		841: note_dur = CYCLES_PER_US * 781;
		842: note_dur = CYCLES_PER_US * 186719;
		843: note_dur = CYCLES_PER_US * 781;
		844: note_dur = CYCLES_PER_US * 186719;
		845: note_dur = CYCLES_PER_US * 781;
		846: note_dur = CYCLES_PER_US * 186719;
		847: note_dur = CYCLES_PER_US * 781;
		848: note_dur = CYCLES_PER_US * 186719;
		849: note_dur = CYCLES_PER_US * 781;
		850: note_dur = CYCLES_PER_US * 186719;
		851: note_dur = CYCLES_PER_US * 781;
		852: note_dur = CYCLES_PER_US * 186719;
		853: note_dur = CYCLES_PER_US * 781;
		854: note_dur = CYCLES_PER_US * 186719;
		855: note_dur = CYCLES_PER_US * 781;
		856: note_dur = CYCLES_PER_US * 186719;
		857: note_dur = CYCLES_PER_US * 781;
		858: note_dur = CYCLES_PER_US * 374219;
		859: note_dur = CYCLES_PER_US * 781;
		860: note_dur = CYCLES_PER_US * 186719;
		861: note_dur = CYCLES_PER_US * 781;
		862: note_dur = CYCLES_PER_US * 92969;
		863: note_dur = CYCLES_PER_US * 781;
		864: note_dur = CYCLES_PER_US * 92969;
		865: note_dur = CYCLES_PER_US * 781;
		866: note_dur = CYCLES_PER_US * 374219;
		867: note_dur = CYCLES_PER_US * 781;
		868: note_dur = CYCLES_PER_US * 1124219;
		869: note_dur = CYCLES_PER_US * 781;
		870: note_dur = CYCLES_PER_US * 92969;
		871: note_dur = CYCLES_PER_US * 781;
		872: note_dur = CYCLES_PER_US * 92969;
		873: note_dur = CYCLES_PER_US * 781;
		874: note_dur = CYCLES_PER_US * 92969;
		875: note_dur = CYCLES_PER_US * 781;
		876: note_dur = CYCLES_PER_US * 92969;
		877: note_dur = CYCLES_PER_US * 781;
		878: note_dur = CYCLES_PER_US * 374219;
		879: note_dur = CYCLES_PER_US * 781;
		880: note_dur = CYCLES_PER_US * 1124219;
		881: note_dur = CYCLES_PER_US * 781;
		882: note_dur = CYCLES_PER_US * 92969;
		883: note_dur = CYCLES_PER_US * 781;
		884: note_dur = CYCLES_PER_US * 92969;
		885: note_dur = CYCLES_PER_US * 781;
		886: note_dur = CYCLES_PER_US * 92969;
		887: note_dur = CYCLES_PER_US * 781;
		888: note_dur = CYCLES_PER_US * 92969;
		889: note_dur = CYCLES_PER_US * 781;
		890: note_dur = CYCLES_PER_US * 374219;
		891: note_dur = CYCLES_PER_US * 781;
		892: note_dur = CYCLES_PER_US * 1124219;
		893: note_dur = CYCLES_PER_US * 1875781;
		894: note_dur = CYCLES_PER_US * 92969;
		895: note_dur = CYCLES_PER_US * 781;
		896: note_dur = CYCLES_PER_US * 92969;
		897: note_dur = CYCLES_PER_US * 781;
		898: note_dur = CYCLES_PER_US * 92969;
		899: note_dur = CYCLES_PER_US * 781;
		900: note_dur = CYCLES_PER_US * 92969;
		901: note_dur = CYCLES_PER_US * 781;
		902: note_dur = CYCLES_PER_US * 374219;
		903: note_dur = CYCLES_PER_US * 781;
		904: note_dur = CYCLES_PER_US * 1124219;
		905: note_dur = CYCLES_PER_US * 1875781;
		906: note_dur = CYCLES_PER_US * 92969;
		907: note_dur = CYCLES_PER_US * 781;
		908: note_dur = CYCLES_PER_US * 92969;
		909: note_dur = CYCLES_PER_US * 781;
		910: note_dur = CYCLES_PER_US * 92969;
		911: note_dur = CYCLES_PER_US * 781;
		912: note_dur = CYCLES_PER_US * 92969;
		913: note_dur = CYCLES_PER_US * 781;
		914: note_dur = CYCLES_PER_US * 374219;
		915: note_dur = CYCLES_PER_US * 781;
		916: note_dur = CYCLES_PER_US * 1124219;
		917: note_dur = CYCLES_PER_US * 1875781;
		918: note_dur = CYCLES_PER_US * 92969;
		919: note_dur = CYCLES_PER_US * 781;
		920: note_dur = CYCLES_PER_US * 92969;
		921: note_dur = CYCLES_PER_US * 781;
		922: note_dur = CYCLES_PER_US * 92969;
		923: note_dur = CYCLES_PER_US * 781;
		924: note_dur = CYCLES_PER_US * 92969;
		925: note_dur = CYCLES_PER_US * 781;
		926: note_dur = CYCLES_PER_US * 374219;
		927: note_dur = CYCLES_PER_US * 0;
		928: note_dur = CYCLES_PER_US * 0;
		929: note_dur = CYCLES_PER_US * 0;
		default: note_dur = 0;
	endcase
end
endmodule