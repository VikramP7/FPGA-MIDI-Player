module song4_dur #(
	parameter int CLOCK_FREQ = 100_000_000
) (
	input logic [10:0] note_index,
	output logic [28:0] note_dur // max 10s at 100MHz clock
);

localparam real TEMPO_BPM = 120;
localparam real CYCLES_PER_BEAT = CLOCK_FREQ*(60/TEMPO_BPM);
localparam real CYCLES_PER_US = CLOCK_FREQ/1000_000;

always_comb begin
	// the quarter note is one beat and therfore can be multipled by CYCLES_PER_BEAT
	case (note_index)
		0: note_dur = CYCLES_PER_US * 416232;
		1: note_dur = CYCLES_PER_US * 434;
		2: note_dur = CYCLES_PER_US * 416232;
		3: note_dur = CYCLES_PER_US * 434;
		4: note_dur = CYCLES_PER_US * 416232;
		5: note_dur = CYCLES_PER_US * 434;
		6: note_dur = CYCLES_PER_US * 312065;
		7: note_dur = CYCLES_PER_US * 434;
		8: note_dur = CYCLES_PER_US * 937064;
		9: note_dur = CYCLES_PER_US * 434;
		10: note_dur = CYCLES_PER_US * 312065;
		11: note_dur = CYCLES_PER_US * 434;
		12: note_dur = CYCLES_PER_US * 520398;
		13: note_dur = CYCLES_PER_US * 434;
		14: note_dur = CYCLES_PER_US * 416232;
		15: note_dur = CYCLES_PER_US * 434;
		16: note_dur = CYCLES_PER_US * 416232;
		17: note_dur = CYCLES_PER_US * 434;
		18: note_dur = CYCLES_PER_US * 416232;
		19: note_dur = CYCLES_PER_US * 434;
		20: note_dur = CYCLES_PER_US * 312065;
		21: note_dur = CYCLES_PER_US * 434;
		22: note_dur = CYCLES_PER_US * 937064;
		23: note_dur = CYCLES_PER_US * 434;
		24: note_dur = CYCLES_PER_US * 416232;
		25: note_dur = CYCLES_PER_US * 434;
		26: note_dur = CYCLES_PER_US * 312065;
		27: note_dur = CYCLES_PER_US * 434;
		28: note_dur = CYCLES_PER_US * 937064;
		29: note_dur = CYCLES_PER_US * 434;
		30: note_dur = CYCLES_PER_US * 416232;
		31: note_dur = CYCLES_PER_US * 434;
		32: note_dur = CYCLES_PER_US * 312065;
		33: note_dur = CYCLES_PER_US * 434;
		34: note_dur = CYCLES_PER_US * 937064;
		35: note_dur = CYCLES_PER_US * 434;
		36: note_dur = CYCLES_PER_US * 416232;
		37: note_dur = CYCLES_PER_US * 434;
		38: note_dur = CYCLES_PER_US * 312065;
		39: note_dur = CYCLES_PER_US * 434;
		40: note_dur = CYCLES_PER_US * 937064;
		41: note_dur = CYCLES_PER_US * 434;
		42: note_dur = CYCLES_PER_US * 416232;
		43: note_dur = CYCLES_PER_US * 434;
		44: note_dur = CYCLES_PER_US * 312065;
		45: note_dur = CYCLES_PER_US * 434;
		46: note_dur = CYCLES_PER_US * 937064;
		47: note_dur = CYCLES_PER_US * 434;
		48: note_dur = CYCLES_PER_US * 312065;
		49: note_dur = CYCLES_PER_US * 434;
		50: note_dur = CYCLES_PER_US * 103732;
		51: note_dur = CYCLES_PER_US * 0;
		52: note_dur = CYCLES_PER_US * 416232;
		53: note_dur = CYCLES_PER_US * 434;
		54: note_dur = CYCLES_PER_US * 416232;
		55: note_dur = CYCLES_PER_US * 434;
		56: note_dur = CYCLES_PER_US * 416232;
		57: note_dur = CYCLES_PER_US * 434;
		58: note_dur = CYCLES_PER_US * 312065;
		59: note_dur = CYCLES_PER_US * 434;
		60: note_dur = CYCLES_PER_US * 937064;
		61: note_dur = CYCLES_PER_US * 434;
		62: note_dur = CYCLES_PER_US * 312065;
		63: note_dur = CYCLES_PER_US * 434;
		64: note_dur = CYCLES_PER_US * 520398;
		65: note_dur = CYCLES_PER_US * 434;
		66: note_dur = CYCLES_PER_US * 416232;
		67: note_dur = CYCLES_PER_US * 434;
		68: note_dur = CYCLES_PER_US * 416232;
		69: note_dur = CYCLES_PER_US * 434;
		70: note_dur = CYCLES_PER_US * 416232;
		71: note_dur = CYCLES_PER_US * 434;
		72: note_dur = CYCLES_PER_US * 312065;
		73: note_dur = CYCLES_PER_US * 434;
		74: note_dur = CYCLES_PER_US * 937064;
		75: note_dur = CYCLES_PER_US * 434;
		76: note_dur = CYCLES_PER_US * 416232;
		77: note_dur = CYCLES_PER_US * 434;
		78: note_dur = CYCLES_PER_US * 312065;
		79: note_dur = CYCLES_PER_US * 434;
		80: note_dur = CYCLES_PER_US * 937064;
		81: note_dur = CYCLES_PER_US * 434;
		82: note_dur = CYCLES_PER_US * 416232;
		83: note_dur = CYCLES_PER_US * 434;
		84: note_dur = CYCLES_PER_US * 312065;
		85: note_dur = CYCLES_PER_US * 434;
		86: note_dur = CYCLES_PER_US * 937064;
		87: note_dur = CYCLES_PER_US * 434;
		88: note_dur = CYCLES_PER_US * 416232;
		89: note_dur = CYCLES_PER_US * 434;
		90: note_dur = CYCLES_PER_US * 312065;
		91: note_dur = CYCLES_PER_US * 434;
		92: note_dur = CYCLES_PER_US * 937064;
		93: note_dur = CYCLES_PER_US * 434;
		94: note_dur = CYCLES_PER_US * 416232;
		95: note_dur = CYCLES_PER_US * 434;
		96: note_dur = CYCLES_PER_US * 312065;
		97: note_dur = CYCLES_PER_US * 434;
		98: note_dur = CYCLES_PER_US * 937064;
		99: note_dur = CYCLES_PER_US * 0;
		100: note_dur = CYCLES_PER_US * 103732;
		101: note_dur = CYCLES_PER_US * 434;
		102: note_dur = CYCLES_PER_US * 103732;
		103: note_dur = CYCLES_PER_US * 434;
		104: note_dur = CYCLES_PER_US * 103732;
		105: note_dur = CYCLES_PER_US * 434;
		106: note_dur = CYCLES_PER_US * 103732;
		107: note_dur = CYCLES_PER_US * 434;
		108: note_dur = CYCLES_PER_US * 312065;
		109: note_dur = CYCLES_PER_US * 434;
		110: note_dur = CYCLES_PER_US * 103732;
		111: note_dur = CYCLES_PER_US * 434;
		112: note_dur = CYCLES_PER_US * 103732;
		113: note_dur = CYCLES_PER_US * 434;
		114: note_dur = CYCLES_PER_US * 103732;
		115: note_dur = CYCLES_PER_US * 434;
		116: note_dur = CYCLES_PER_US * 207899;
		117: note_dur = CYCLES_PER_US * 434;
		118: note_dur = CYCLES_PER_US * 103732;
		119: note_dur = CYCLES_PER_US * 434;
		120: note_dur = CYCLES_PER_US * 103732;
		121: note_dur = CYCLES_PER_US * 434;
		122: note_dur = CYCLES_PER_US * 103732;
		123: note_dur = CYCLES_PER_US * 434;
		124: note_dur = CYCLES_PER_US * 103732;
		125: note_dur = CYCLES_PER_US * 434;
		126: note_dur = CYCLES_PER_US * 103732;
		127: note_dur = CYCLES_PER_US * 434;
		128: note_dur = CYCLES_PER_US * 103732;
		129: note_dur = CYCLES_PER_US * 434;
		130: note_dur = CYCLES_PER_US * 207899;
		131: note_dur = CYCLES_PER_US * 434;
		132: note_dur = CYCLES_PER_US * 103732;
		133: note_dur = CYCLES_PER_US * 434;
		134: note_dur = CYCLES_PER_US * 103732;
		135: note_dur = CYCLES_PER_US * 434;
		136: note_dur = CYCLES_PER_US * 103732;
		137: note_dur = CYCLES_PER_US * 434;
		138: note_dur = CYCLES_PER_US * 103732;
		139: note_dur = CYCLES_PER_US * 434;
		140: note_dur = CYCLES_PER_US * 103732;
		141: note_dur = CYCLES_PER_US * 434;
		142: note_dur = CYCLES_PER_US * 103732;
		143: note_dur = CYCLES_PER_US * 434;
		144: note_dur = CYCLES_PER_US * 103732;
		145: note_dur = CYCLES_PER_US * 434;
		146: note_dur = CYCLES_PER_US * 103732;
		147: note_dur = CYCLES_PER_US * 434;
		148: note_dur = CYCLES_PER_US * 103732;
		149: note_dur = CYCLES_PER_US * 434;
		150: note_dur = CYCLES_PER_US * 103732;
		151: note_dur = CYCLES_PER_US * 434;
		152: note_dur = CYCLES_PER_US * 103732;
		153: note_dur = CYCLES_PER_US * 434;
		154: note_dur = CYCLES_PER_US * 103732;
		155: note_dur = CYCLES_PER_US * 434;
		156: note_dur = CYCLES_PER_US * 103732;
		157: note_dur = CYCLES_PER_US * 434;
		158: note_dur = CYCLES_PER_US * 103732;
		159: note_dur = CYCLES_PER_US * 434;
		160: note_dur = CYCLES_PER_US * 103732;
		161: note_dur = CYCLES_PER_US * 434;
		162: note_dur = CYCLES_PER_US * 103732;
		163: note_dur = CYCLES_PER_US * 434;
		164: note_dur = CYCLES_PER_US * 103732;
		165: note_dur = CYCLES_PER_US * 434;
		166: note_dur = CYCLES_PER_US * 103732;
		167: note_dur = CYCLES_PER_US * 434;
		168: note_dur = CYCLES_PER_US * 103732;
		169: note_dur = CYCLES_PER_US * 434;
		170: note_dur = CYCLES_PER_US * 103732;
		171: note_dur = CYCLES_PER_US * 434;
		172: note_dur = CYCLES_PER_US * 103732;
		173: note_dur = CYCLES_PER_US * 434;
		174: note_dur = CYCLES_PER_US * 103732;
		175: note_dur = CYCLES_PER_US * 434;
		176: note_dur = CYCLES_PER_US * 103732;
		177: note_dur = CYCLES_PER_US * 434;
		178: note_dur = CYCLES_PER_US * 103732;
		179: note_dur = CYCLES_PER_US * 434;
		180: note_dur = CYCLES_PER_US * 103732;
		181: note_dur = CYCLES_PER_US * 434;
		182: note_dur = CYCLES_PER_US * 103732;
		183: note_dur = CYCLES_PER_US * 434;
		184: note_dur = CYCLES_PER_US * 103732;
		185: note_dur = CYCLES_PER_US * 434;
		186: note_dur = CYCLES_PER_US * 103732;
		187: note_dur = CYCLES_PER_US * 434;
		188: note_dur = CYCLES_PER_US * 103732;
		189: note_dur = CYCLES_PER_US * 434;
		190: note_dur = CYCLES_PER_US * 103732;
		191: note_dur = CYCLES_PER_US * 434;
		192: note_dur = CYCLES_PER_US * 103732;
		193: note_dur = CYCLES_PER_US * 434;
		194: note_dur = CYCLES_PER_US * 103732;
		195: note_dur = CYCLES_PER_US * 434;
		196: note_dur = CYCLES_PER_US * 103732;
		197: note_dur = CYCLES_PER_US * 434;
		198: note_dur = CYCLES_PER_US * 103732;
		199: note_dur = CYCLES_PER_US * 434;
		200: note_dur = CYCLES_PER_US * 103732;
		201: note_dur = CYCLES_PER_US * 434;
		202: note_dur = CYCLES_PER_US * 103732;
		203: note_dur = CYCLES_PER_US * 434;
		204: note_dur = CYCLES_PER_US * 207899;
		205: note_dur = CYCLES_PER_US * 434;
		206: note_dur = CYCLES_PER_US * 103732;
		207: note_dur = CYCLES_PER_US * 434;
		208: note_dur = CYCLES_PER_US * 103732;
		209: note_dur = CYCLES_PER_US * 417100;
		210: note_dur = CYCLES_PER_US * 103732;
		211: note_dur = CYCLES_PER_US * 434;
		212: note_dur = CYCLES_PER_US * 103732;
		213: note_dur = CYCLES_PER_US * 434;
		214: note_dur = CYCLES_PER_US * 103732;
		215: note_dur = CYCLES_PER_US * 434;
		216: note_dur = CYCLES_PER_US * 103732;
		217: note_dur = CYCLES_PER_US * 434;
		218: note_dur = CYCLES_PER_US * 103732;
		219: note_dur = CYCLES_PER_US * 434;
		220: note_dur = CYCLES_PER_US * 103732;
		221: note_dur = CYCLES_PER_US * 434;
		222: note_dur = CYCLES_PER_US * 103732;
		223: note_dur = CYCLES_PER_US * 434;
		224: note_dur = CYCLES_PER_US * 103732;
		225: note_dur = CYCLES_PER_US * 434;
		226: note_dur = CYCLES_PER_US * 103732;
		227: note_dur = CYCLES_PER_US * 434;
		228: note_dur = CYCLES_PER_US * 103732;
		229: note_dur = CYCLES_PER_US * 434;
		230: note_dur = CYCLES_PER_US * 103732;
		231: note_dur = CYCLES_PER_US * 434;
		232: note_dur = CYCLES_PER_US * 103732;
		233: note_dur = CYCLES_PER_US * 434;
		234: note_dur = CYCLES_PER_US * 103732;
		235: note_dur = CYCLES_PER_US * 434;
		236: note_dur = CYCLES_PER_US * 103732;
		237: note_dur = CYCLES_PER_US * 434;
		238: note_dur = CYCLES_PER_US * 103732;
		239: note_dur = CYCLES_PER_US * 434;
		240: note_dur = CYCLES_PER_US * 103732;
		241: note_dur = CYCLES_PER_US * 434;
		242: note_dur = CYCLES_PER_US * 103732;
		243: note_dur = CYCLES_PER_US * 434;
		244: note_dur = CYCLES_PER_US * 103732;
		245: note_dur = CYCLES_PER_US * 434;
		246: note_dur = CYCLES_PER_US * 103732;
		247: note_dur = CYCLES_PER_US * 434;
		248: note_dur = CYCLES_PER_US * 103732;
		249: note_dur = CYCLES_PER_US * 434;
		250: note_dur = CYCLES_PER_US * 103732;
		251: note_dur = CYCLES_PER_US * 434;
		252: note_dur = CYCLES_PER_US * 103732;
		253: note_dur = CYCLES_PER_US * 434;
		254: note_dur = CYCLES_PER_US * 103732;
		255: note_dur = CYCLES_PER_US * 434;
		256: note_dur = CYCLES_PER_US * 103732;
		257: note_dur = CYCLES_PER_US * 434;
		258: note_dur = CYCLES_PER_US * 103732;
		259: note_dur = CYCLES_PER_US * 434;
		260: note_dur = CYCLES_PER_US * 103732;
		261: note_dur = CYCLES_PER_US * 434;
		262: note_dur = CYCLES_PER_US * 103732;
		263: note_dur = CYCLES_PER_US * 434;
		264: note_dur = CYCLES_PER_US * 103732;
		265: note_dur = CYCLES_PER_US * 434;
		266: note_dur = CYCLES_PER_US * 103732;
		267: note_dur = CYCLES_PER_US * 434;
		268: note_dur = CYCLES_PER_US * 103732;
		269: note_dur = CYCLES_PER_US * 434;
		270: note_dur = CYCLES_PER_US * 103732;
		271: note_dur = CYCLES_PER_US * 434;
		272: note_dur = CYCLES_PER_US * 103732;
		273: note_dur = CYCLES_PER_US * 434;
		274: note_dur = CYCLES_PER_US * 103732;
		275: note_dur = CYCLES_PER_US * 434;
		276: note_dur = CYCLES_PER_US * 103732;
		277: note_dur = CYCLES_PER_US * 434;
		278: note_dur = CYCLES_PER_US * 103732;
		279: note_dur = CYCLES_PER_US * 434;
		280: note_dur = CYCLES_PER_US * 207899;
		281: note_dur = CYCLES_PER_US * 434;
		282: note_dur = CYCLES_PER_US * 103732;
		283: note_dur = CYCLES_PER_US * 434;
		284: note_dur = CYCLES_PER_US * 103732;
		285: note_dur = CYCLES_PER_US * 434;
		286: note_dur = CYCLES_PER_US * 103732;
		287: note_dur = CYCLES_PER_US * 434;
		288: note_dur = CYCLES_PER_US * 103732;
		289: note_dur = CYCLES_PER_US * 434;
		290: note_dur = CYCLES_PER_US * 103732;
		291: note_dur = CYCLES_PER_US * 434;
		292: note_dur = CYCLES_PER_US * 103732;
		293: note_dur = CYCLES_PER_US * 434;
		294: note_dur = CYCLES_PER_US * 103732;
		295: note_dur = CYCLES_PER_US * 434;
		296: note_dur = CYCLES_PER_US * 103732;
		297: note_dur = CYCLES_PER_US * 434;
		298: note_dur = CYCLES_PER_US * 103732;
		299: note_dur = CYCLES_PER_US * 434;
		300: note_dur = CYCLES_PER_US * 103732;
		301: note_dur = CYCLES_PER_US * 434;
		302: note_dur = CYCLES_PER_US * 103732;
		303: note_dur = CYCLES_PER_US * 434;
		304: note_dur = CYCLES_PER_US * 207899;
		305: note_dur = CYCLES_PER_US * 208767;
		306: note_dur = CYCLES_PER_US * 103732;
		307: note_dur = CYCLES_PER_US * 434;
		308: note_dur = CYCLES_PER_US * 103732;
		309: note_dur = CYCLES_PER_US * 434;
		310: note_dur = CYCLES_PER_US * 103732;
		311: note_dur = CYCLES_PER_US * 434;
		312: note_dur = CYCLES_PER_US * 103732;
		313: note_dur = CYCLES_PER_US * 434;
		314: note_dur = CYCLES_PER_US * 103732;
		315: note_dur = CYCLES_PER_US * 434;
		316: note_dur = CYCLES_PER_US * 103732;
		317: note_dur = CYCLES_PER_US * 434;
		318: note_dur = CYCLES_PER_US * 103732;
		319: note_dur = CYCLES_PER_US * 434;
		320: note_dur = CYCLES_PER_US * 103732;
		321: note_dur = CYCLES_PER_US * 434;
		322: note_dur = CYCLES_PER_US * 103732;
		323: note_dur = CYCLES_PER_US * 434;
		324: note_dur = CYCLES_PER_US * 103732;
		325: note_dur = CYCLES_PER_US * 486544;
		326: note_dur = CYCLES_PER_US * 69010;
		327: note_dur = CYCLES_PER_US * 434;
		328: note_dur = CYCLES_PER_US * 69010;
		329: note_dur = CYCLES_PER_US * 434;
		330: note_dur = CYCLES_PER_US * 312065;
		331: note_dur = CYCLES_PER_US * 434;
		332: note_dur = CYCLES_PER_US * 103732;
		333: note_dur = CYCLES_PER_US * 434;
		334: note_dur = CYCLES_PER_US * 0;
		335: note_dur = CYCLES_PER_US * 0;
		336: note_dur = CYCLES_PER_US * 0;
		337: note_dur = CYCLES_PER_US * 624565;
		338: note_dur = CYCLES_PER_US * 0;
		339: note_dur = CYCLES_PER_US * 0;
		340: note_dur = CYCLES_PER_US * 0;
		341: note_dur = CYCLES_PER_US * 104601;
		342: note_dur = CYCLES_PER_US * 103732;
		343: note_dur = CYCLES_PER_US * 434;
		344: note_dur = CYCLES_PER_US * 103732;
		345: note_dur = CYCLES_PER_US * 434;
		346: note_dur = CYCLES_PER_US * 103732;
		347: note_dur = CYCLES_PER_US * 434;
		348: note_dur = CYCLES_PER_US * 103732;
		349: note_dur = CYCLES_PER_US * 434;
		350: note_dur = CYCLES_PER_US * 103732;
		351: note_dur = CYCLES_PER_US * 434;
		352: note_dur = CYCLES_PER_US * 103732;
		353: note_dur = CYCLES_PER_US * 434;
		354: note_dur = CYCLES_PER_US * 103732;
		355: note_dur = CYCLES_PER_US * 434;
		356: note_dur = CYCLES_PER_US * 103732;
		357: note_dur = CYCLES_PER_US * 434;
		358: note_dur = CYCLES_PER_US * 103732;
		359: note_dur = CYCLES_PER_US * 434;
		360: note_dur = CYCLES_PER_US * 103732;
		361: note_dur = CYCLES_PER_US * 434;
		362: note_dur = CYCLES_PER_US * 103732;
		363: note_dur = CYCLES_PER_US * 434;
		364: note_dur = CYCLES_PER_US * 103732;
		365: note_dur = CYCLES_PER_US * 434;
		366: note_dur = CYCLES_PER_US * 103732;
		367: note_dur = CYCLES_PER_US * 434;
		368: note_dur = CYCLES_PER_US * 103732;
		369: note_dur = CYCLES_PER_US * 434;
		370: note_dur = CYCLES_PER_US * 103732;
		371: note_dur = CYCLES_PER_US * 208767;
		372: note_dur = CYCLES_PER_US * 0;
		373: note_dur = CYCLES_PER_US * 0;
		374: note_dur = CYCLES_PER_US * 0;
		375: note_dur = CYCLES_PER_US * 0;
		376: note_dur = CYCLES_PER_US * 312065;
		377: note_dur = CYCLES_PER_US * 0;
		378: note_dur = CYCLES_PER_US * 0;
		379: note_dur = CYCLES_PER_US * 0;
		380: note_dur = CYCLES_PER_US * 0;
		381: note_dur = CYCLES_PER_US * 434;
		382: note_dur = CYCLES_PER_US * 207899;
		383: note_dur = CYCLES_PER_US * 434;
		384: note_dur = CYCLES_PER_US * 103732;
		385: note_dur = CYCLES_PER_US * 434;
		386: note_dur = CYCLES_PER_US * 207899;
		387: note_dur = CYCLES_PER_US * 104601;
		388: note_dur = CYCLES_PER_US * 103732;
		389: note_dur = CYCLES_PER_US * 434;
		390: note_dur = CYCLES_PER_US * 103732;
		391: note_dur = CYCLES_PER_US * 434;
		392: note_dur = CYCLES_PER_US * 103732;
		393: note_dur = CYCLES_PER_US * 434;
		394: note_dur = CYCLES_PER_US * 103732;
		395: note_dur = CYCLES_PER_US * 434;
		396: note_dur = CYCLES_PER_US * 103732;
		397: note_dur = CYCLES_PER_US * 434;
		398: note_dur = CYCLES_PER_US * 103732;
		399: note_dur = CYCLES_PER_US * 434;
		400: note_dur = CYCLES_PER_US * 103732;
		401: note_dur = CYCLES_PER_US * 434;
		402: note_dur = CYCLES_PER_US * 103732;
		403: note_dur = CYCLES_PER_US * 434;
		404: note_dur = CYCLES_PER_US * 103732;
		405: note_dur = CYCLES_PER_US * 434;
		406: note_dur = CYCLES_PER_US * 103732;
		407: note_dur = CYCLES_PER_US * 434;
		408: note_dur = CYCLES_PER_US * 103732;
		409: note_dur = CYCLES_PER_US * 434;
		410: note_dur = CYCLES_PER_US * 103732;
		411: note_dur = CYCLES_PER_US * 434;
		412: note_dur = CYCLES_PER_US * 103732;
		413: note_dur = CYCLES_PER_US * 434;
		414: note_dur = CYCLES_PER_US * 103732;
		415: note_dur = CYCLES_PER_US * 434;
		416: note_dur = CYCLES_PER_US * 103732;
		417: note_dur = CYCLES_PER_US * 434;
		418: note_dur = CYCLES_PER_US * 312065;
		419: note_dur = CYCLES_PER_US * 434;
		420: note_dur = CYCLES_PER_US * 103732;
		421: note_dur = CYCLES_PER_US * 434;
		422: note_dur = CYCLES_PER_US * 103732;
		423: note_dur = CYCLES_PER_US * 434;
		424: note_dur = CYCLES_PER_US * 103732;
		425: note_dur = CYCLES_PER_US * 434;
		426: note_dur = CYCLES_PER_US * 103732;
		427: note_dur = CYCLES_PER_US * 434;
		428: note_dur = CYCLES_PER_US * 103732;
		429: note_dur = CYCLES_PER_US * 434;
		430: note_dur = CYCLES_PER_US * 103732;
		431: note_dur = CYCLES_PER_US * 434;
		432: note_dur = CYCLES_PER_US * 103732;
		433: note_dur = CYCLES_PER_US * 434;
		434: note_dur = CYCLES_PER_US * 103732;
		435: note_dur = CYCLES_PER_US * 434;
		436: note_dur = CYCLES_PER_US * 103732;
		437: note_dur = CYCLES_PER_US * 434;
		438: note_dur = CYCLES_PER_US * 103732;
		439: note_dur = CYCLES_PER_US * 434;
		440: note_dur = CYCLES_PER_US * 103732;
		441: note_dur = CYCLES_PER_US * 434;
		442: note_dur = CYCLES_PER_US * 103732;
		443: note_dur = CYCLES_PER_US * 434;
		444: note_dur = CYCLES_PER_US * 103732;
		445: note_dur = CYCLES_PER_US * 434;
		446: note_dur = CYCLES_PER_US * 207899;
		447: note_dur = CYCLES_PER_US * 104601;
		448: note_dur = CYCLES_PER_US * 103732;
		449: note_dur = CYCLES_PER_US * 434;
		450: note_dur = CYCLES_PER_US * 103732;
		451: note_dur = CYCLES_PER_US * 434;
		452: note_dur = CYCLES_PER_US * 103732;
		453: note_dur = CYCLES_PER_US * 312934;
		454: note_dur = CYCLES_PER_US * 103732;
		455: note_dur = CYCLES_PER_US * 434;
		456: note_dur = CYCLES_PER_US * 103732;
		457: note_dur = CYCLES_PER_US * 434;
		458: note_dur = CYCLES_PER_US * 103732;
		459: note_dur = CYCLES_PER_US * 434;
		460: note_dur = CYCLES_PER_US * 103732;
		461: note_dur = CYCLES_PER_US * 434;
		462: note_dur = CYCLES_PER_US * 103732;
		463: note_dur = CYCLES_PER_US * 434;
		464: note_dur = CYCLES_PER_US * 103732;
		465: note_dur = CYCLES_PER_US * 434;
		466: note_dur = CYCLES_PER_US * 103732;
		467: note_dur = CYCLES_PER_US * 434;
		468: note_dur = CYCLES_PER_US * 103732;
		469: note_dur = CYCLES_PER_US * 434;
		470: note_dur = CYCLES_PER_US * 103732;
		471: note_dur = CYCLES_PER_US * 434;
		472: note_dur = CYCLES_PER_US * 103732;
		473: note_dur = CYCLES_PER_US * 434;
		474: note_dur = CYCLES_PER_US * 103732;
		475: note_dur = CYCLES_PER_US * 434;
		476: note_dur = CYCLES_PER_US * 103732;
		477: note_dur = CYCLES_PER_US * 434;
		478: note_dur = CYCLES_PER_US * 103732;
		479: note_dur = CYCLES_PER_US * 434;
		480: note_dur = CYCLES_PER_US * 103732;
		481: note_dur = CYCLES_PER_US * 434;
		482: note_dur = CYCLES_PER_US * 207899;
		483: note_dur = CYCLES_PER_US * 434;
		484: note_dur = CYCLES_PER_US * 416232;
		485: note_dur = CYCLES_PER_US * 312934;
		486: note_dur = CYCLES_PER_US * 103732;
		487: note_dur = CYCLES_PER_US * 434;
		488: note_dur = CYCLES_PER_US * 103732;
		489: note_dur = CYCLES_PER_US * 434;
		490: note_dur = CYCLES_PER_US * 103732;
		491: note_dur = CYCLES_PER_US * 434;
		492: note_dur = CYCLES_PER_US * 103732;
		493: note_dur = CYCLES_PER_US * 434;
		494: note_dur = CYCLES_PER_US * 103732;
		495: note_dur = CYCLES_PER_US * 434;
		496: note_dur = CYCLES_PER_US * 103732;
		497: note_dur = CYCLES_PER_US * 434;
		498: note_dur = CYCLES_PER_US * 103732;
		499: note_dur = CYCLES_PER_US * 434;
		500: note_dur = CYCLES_PER_US * 103732;
		501: note_dur = CYCLES_PER_US * 434;
		502: note_dur = CYCLES_PER_US * 103732;
		503: note_dur = CYCLES_PER_US * 434;
		504: note_dur = CYCLES_PER_US * 103732;
		505: note_dur = CYCLES_PER_US * 434;
		506: note_dur = CYCLES_PER_US * 103732;
		507: note_dur = CYCLES_PER_US * 434;
		508: note_dur = CYCLES_PER_US * 103732;
		509: note_dur = CYCLES_PER_US * 434;
		510: note_dur = CYCLES_PER_US * 103732;
		511: note_dur = CYCLES_PER_US * 434;
		512: note_dur = CYCLES_PER_US * 103732;
		513: note_dur = CYCLES_PER_US * 434;
		514: note_dur = CYCLES_PER_US * 103732;
		515: note_dur = CYCLES_PER_US * 434;
		516: note_dur = CYCLES_PER_US * 103732;
		517: note_dur = CYCLES_PER_US * 434;
		518: note_dur = CYCLES_PER_US * 312065;
		519: note_dur = CYCLES_PER_US * 434;
		520: note_dur = CYCLES_PER_US * 312065;
		521: note_dur = CYCLES_PER_US * 312934;
		522: note_dur = CYCLES_PER_US * 103732;
		523: note_dur = CYCLES_PER_US * 434;
		524: note_dur = CYCLES_PER_US * 69010;
		525: note_dur = CYCLES_PER_US * 434;
		526: note_dur = CYCLES_PER_US * 69010;
		527: note_dur = CYCLES_PER_US * 434;
		528: note_dur = CYCLES_PER_US * 69010;
		529: note_dur = CYCLES_PER_US * 434;
		530: note_dur = CYCLES_PER_US * 103732;
		531: note_dur = CYCLES_PER_US * 434;
		532: note_dur = CYCLES_PER_US * 103732;
		533: note_dur = CYCLES_PER_US * 434;
		534: note_dur = CYCLES_PER_US * 103732;
		535: note_dur = CYCLES_PER_US * 434;
		536: note_dur = CYCLES_PER_US * 103732;
		537: note_dur = CYCLES_PER_US * 434;
		538: note_dur = CYCLES_PER_US * 0;
		539: note_dur = CYCLES_PER_US * 103732;
		540: note_dur = CYCLES_PER_US * 0;
		541: note_dur = CYCLES_PER_US * 434;
		542: note_dur = CYCLES_PER_US * 103732;
		543: note_dur = CYCLES_PER_US * 434;
		544: note_dur = CYCLES_PER_US * 103732;
		545: note_dur = CYCLES_PER_US * 434;
		546: note_dur = CYCLES_PER_US * 103732;
		547: note_dur = CYCLES_PER_US * 434;
		548: note_dur = CYCLES_PER_US * 103732;
		549: note_dur = CYCLES_PER_US * 434;
		550: note_dur = CYCLES_PER_US * 103732;
		551: note_dur = CYCLES_PER_US * 434;
		552: note_dur = CYCLES_PER_US * 103732;
		553: note_dur = CYCLES_PER_US * 434;
		554: note_dur = CYCLES_PER_US * 103732;
		555: note_dur = CYCLES_PER_US * 434;
		556: note_dur = CYCLES_PER_US * 103732;
		557: note_dur = CYCLES_PER_US * 434;
		558: note_dur = CYCLES_PER_US * 103732;
		559: note_dur = CYCLES_PER_US * 434;
		560: note_dur = CYCLES_PER_US * 207899;
		561: note_dur = CYCLES_PER_US * 434;
		562: note_dur = CYCLES_PER_US * 103732;
		563: note_dur = CYCLES_PER_US * 434;
		564: note_dur = CYCLES_PER_US * 103732;
		565: note_dur = CYCLES_PER_US * 434;
		566: note_dur = CYCLES_PER_US * 103732;
		567: note_dur = CYCLES_PER_US * 434;
		568: note_dur = CYCLES_PER_US * 103732;
		569: note_dur = CYCLES_PER_US * 434;
		570: note_dur = CYCLES_PER_US * 103732;
		571: note_dur = CYCLES_PER_US * 434;
		572: note_dur = CYCLES_PER_US * 103732;
		573: note_dur = CYCLES_PER_US * 434;
		574: note_dur = CYCLES_PER_US * 103732;
		575: note_dur = CYCLES_PER_US * 434;
		576: note_dur = CYCLES_PER_US * 103732;
		577: note_dur = CYCLES_PER_US * 434;
		578: note_dur = CYCLES_PER_US * 103732;
		579: note_dur = CYCLES_PER_US * 434;
		580: note_dur = CYCLES_PER_US * 103732;
		581: note_dur = CYCLES_PER_US * 434;
		582: note_dur = CYCLES_PER_US * 103732;
		583: note_dur = CYCLES_PER_US * 434;
		584: note_dur = CYCLES_PER_US * 103732;
		585: note_dur = CYCLES_PER_US * 434;
		586: note_dur = CYCLES_PER_US * 103732;
		587: note_dur = CYCLES_PER_US * 434;
		588: note_dur = CYCLES_PER_US * 103732;
		589: note_dur = CYCLES_PER_US * 208767;
		590: note_dur = CYCLES_PER_US * 103732;
		591: note_dur = CYCLES_PER_US * 434;
		592: note_dur = CYCLES_PER_US * 103732;
		593: note_dur = CYCLES_PER_US * 434;
		594: note_dur = CYCLES_PER_US * 103732;
		595: note_dur = CYCLES_PER_US * 434;
		596: note_dur = CYCLES_PER_US * 103732;
		597: note_dur = CYCLES_PER_US * 434;
		598: note_dur = CYCLES_PER_US * 103732;
		599: note_dur = CYCLES_PER_US * 434;
		600: note_dur = CYCLES_PER_US * 103732;
		601: note_dur = CYCLES_PER_US * 434;
		602: note_dur = CYCLES_PER_US * 103732;
		603: note_dur = CYCLES_PER_US * 434;
		604: note_dur = CYCLES_PER_US * 103732;
		605: note_dur = CYCLES_PER_US * 434;
		606: note_dur = CYCLES_PER_US * 103732;
		607: note_dur = CYCLES_PER_US * 434;
		608: note_dur = CYCLES_PER_US * 103732;
		609: note_dur = CYCLES_PER_US * 434;
		610: note_dur = CYCLES_PER_US * 103732;
		611: note_dur = CYCLES_PER_US * 434;
		612: note_dur = CYCLES_PER_US * 103732;
		613: note_dur = CYCLES_PER_US * 434;
		614: note_dur = CYCLES_PER_US * 103732;
		615: note_dur = CYCLES_PER_US * 434;
		616: note_dur = CYCLES_PER_US * 103732;
		617: note_dur = CYCLES_PER_US * 434;
		618: note_dur = CYCLES_PER_US * 103732;
		619: note_dur = CYCLES_PER_US * 434;
		620: note_dur = CYCLES_PER_US * 103732;
		621: note_dur = CYCLES_PER_US * 434;
		622: note_dur = CYCLES_PER_US * 103732;
		623: note_dur = CYCLES_PER_US * 434;
		624: note_dur = CYCLES_PER_US * 103732;
		625: note_dur = CYCLES_PER_US * 434;
		626: note_dur = CYCLES_PER_US * 103732;
		627: note_dur = CYCLES_PER_US * 434;
		628: note_dur = CYCLES_PER_US * 103732;
		629: note_dur = CYCLES_PER_US * 434;
		630: note_dur = CYCLES_PER_US * 207899;
		631: note_dur = CYCLES_PER_US * 434;
		632: note_dur = CYCLES_PER_US * 103732;
		633: note_dur = CYCLES_PER_US * 434;
		634: note_dur = CYCLES_PER_US * 103732;
		635: note_dur = CYCLES_PER_US * 434;
		636: note_dur = CYCLES_PER_US * 103732;
		637: note_dur = CYCLES_PER_US * 434;
		638: note_dur = CYCLES_PER_US * 103732;
		639: note_dur = CYCLES_PER_US * 521267;
		640: note_dur = CYCLES_PER_US * 0;
		641: note_dur = CYCLES_PER_US * 0;
		642: note_dur = CYCLES_PER_US * 0;
		643: note_dur = CYCLES_PER_US * 0;
		644: note_dur = CYCLES_PER_US * 103732;
		645: note_dur = CYCLES_PER_US * 0;
		646: note_dur = CYCLES_PER_US * 0;
		647: note_dur = CYCLES_PER_US * 0;
		648: note_dur = CYCLES_PER_US * 312500;
		649: note_dur = CYCLES_PER_US * 434;
		650: note_dur = CYCLES_PER_US * 51649;
		651: note_dur = CYCLES_PER_US * 434;
		652: note_dur = CYCLES_PER_US * 51649;
		653: note_dur = CYCLES_PER_US * 434;
		654: note_dur = CYCLES_PER_US * 103732;
		655: note_dur = CYCLES_PER_US * 434;
		656: note_dur = CYCLES_PER_US * 103732;
		657: note_dur = CYCLES_PER_US * 434;
		658: note_dur = CYCLES_PER_US * 103732;
		659: note_dur = CYCLES_PER_US * 434;
		660: note_dur = CYCLES_PER_US * 103732;
		661: note_dur = CYCLES_PER_US * 434;
		662: note_dur = CYCLES_PER_US * 103732;
		663: note_dur = CYCLES_PER_US * 434;
		664: note_dur = CYCLES_PER_US * 103732;
		665: note_dur = CYCLES_PER_US * 434;
		666: note_dur = CYCLES_PER_US * 103732;
		667: note_dur = CYCLES_PER_US * 434;
		668: note_dur = CYCLES_PER_US * 103732;
		669: note_dur = CYCLES_PER_US * 434;
		670: note_dur = CYCLES_PER_US * 0;
		671: note_dur = CYCLES_PER_US * 0;
		672: note_dur = CYCLES_PER_US * 0;
		673: note_dur = CYCLES_PER_US * 624565;
		674: note_dur = CYCLES_PER_US * 0;
		675: note_dur = CYCLES_PER_US * 0;
		676: note_dur = CYCLES_PER_US * 104166;
		677: note_dur = CYCLES_PER_US * 434;
		678: note_dur = CYCLES_PER_US * 34288;
		679: note_dur = CYCLES_PER_US * 434;
		680: note_dur = CYCLES_PER_US * 34288;
		681: note_dur = CYCLES_PER_US * 434;
		682: note_dur = CYCLES_PER_US * 34288;
		683: note_dur = CYCLES_PER_US * 434;
		684: note_dur = CYCLES_PER_US * 103732;
		685: note_dur = CYCLES_PER_US * 434;
		686: note_dur = CYCLES_PER_US * 103732;
		687: note_dur = CYCLES_PER_US * 434;
		688: note_dur = CYCLES_PER_US * 103732;
		689: note_dur = CYCLES_PER_US * 434;
		690: note_dur = CYCLES_PER_US * 103732;
		691: note_dur = CYCLES_PER_US * 434;
		692: note_dur = CYCLES_PER_US * 103732;
		693: note_dur = CYCLES_PER_US * 434;
		694: note_dur = CYCLES_PER_US * 103732;
		695: note_dur = CYCLES_PER_US * 434;
		696: note_dur = CYCLES_PER_US * 103732;
		697: note_dur = CYCLES_PER_US * 434;
		698: note_dur = CYCLES_PER_US * 103732;
		699: note_dur = CYCLES_PER_US * 434;
		700: note_dur = CYCLES_PER_US * 103732;
		701: note_dur = CYCLES_PER_US * 434;
		702: note_dur = CYCLES_PER_US * 103732;
		703: note_dur = CYCLES_PER_US * 434;
		704: note_dur = CYCLES_PER_US * 103732;
		705: note_dur = CYCLES_PER_US * 434;
		706: note_dur = CYCLES_PER_US * 103732;
		707: note_dur = CYCLES_PER_US * 434;
		708: note_dur = CYCLES_PER_US * 103732;
		709: note_dur = CYCLES_PER_US * 434;
		710: note_dur = CYCLES_PER_US * 103732;
		711: note_dur = CYCLES_PER_US * 434;
		712: note_dur = CYCLES_PER_US * 103732;
		713: note_dur = CYCLES_PER_US * 434;
		714: note_dur = CYCLES_PER_US * 103732;
		715: note_dur = CYCLES_PER_US * 434;
		716: note_dur = CYCLES_PER_US * 103732;
		717: note_dur = CYCLES_PER_US * 434;
		718: note_dur = CYCLES_PER_US * 103732;
		719: note_dur = CYCLES_PER_US * 434;
		720: note_dur = CYCLES_PER_US * 103732;
		721: note_dur = CYCLES_PER_US * 434;
		722: note_dur = CYCLES_PER_US * 103732;
		723: note_dur = CYCLES_PER_US * 434;
		724: note_dur = CYCLES_PER_US * 103732;
		725: note_dur = CYCLES_PER_US * 434;
		726: note_dur = CYCLES_PER_US * 103732;
		727: note_dur = CYCLES_PER_US * 434;
		728: note_dur = CYCLES_PER_US * 103732;
		729: note_dur = CYCLES_PER_US * 434;
		730: note_dur = CYCLES_PER_US * 103732;
		731: note_dur = CYCLES_PER_US * 434;
		732: note_dur = CYCLES_PER_US * 312065;
		733: note_dur = CYCLES_PER_US * 434;
		734: note_dur = CYCLES_PER_US * 51649;
		735: note_dur = CYCLES_PER_US * 434;
		736: note_dur = CYCLES_PER_US * 51649;
		737: note_dur = CYCLES_PER_US * 434;
		738: note_dur = CYCLES_PER_US * 103732;
		739: note_dur = CYCLES_PER_US * 434;
		740: note_dur = CYCLES_PER_US * 103732;
		741: note_dur = CYCLES_PER_US * 434;
		742: note_dur = CYCLES_PER_US * 103732;
		743: note_dur = CYCLES_PER_US * 434;
		744: note_dur = CYCLES_PER_US * 103732;
		745: note_dur = CYCLES_PER_US * 434;
		746: note_dur = CYCLES_PER_US * 103732;
		747: note_dur = CYCLES_PER_US * 434;
		748: note_dur = CYCLES_PER_US * 103732;
		749: note_dur = CYCLES_PER_US * 434;
		750: note_dur = CYCLES_PER_US * 103732;
		751: note_dur = CYCLES_PER_US * 434;
		752: note_dur = CYCLES_PER_US * 103732;
		753: note_dur = CYCLES_PER_US * 434;
		754: note_dur = CYCLES_PER_US * 103732;
		755: note_dur = CYCLES_PER_US * 434;
		756: note_dur = CYCLES_PER_US * 103732;
		757: note_dur = CYCLES_PER_US * 434;
		758: note_dur = CYCLES_PER_US * 103732;
		759: note_dur = CYCLES_PER_US * 434;
		760: note_dur = CYCLES_PER_US * 103732;
		761: note_dur = CYCLES_PER_US * 434;
		762: note_dur = CYCLES_PER_US * 207899;
		763: note_dur = CYCLES_PER_US * 729600;
		764: note_dur = CYCLES_PER_US * 103732;
		765: note_dur = CYCLES_PER_US * 434;
		766: note_dur = CYCLES_PER_US * 103732;
		767: note_dur = CYCLES_PER_US * 434;
		768: note_dur = CYCLES_PER_US * 103732;
		769: note_dur = CYCLES_PER_US * 434;
		770: note_dur = CYCLES_PER_US * 103732;
		771: note_dur = CYCLES_PER_US * 434;
		772: note_dur = CYCLES_PER_US * 103732;
		773: note_dur = CYCLES_PER_US * 434;
		774: note_dur = CYCLES_PER_US * 103732;
		775: note_dur = CYCLES_PER_US * 434;
		776: note_dur = CYCLES_PER_US * 103732;
		777: note_dur = CYCLES_PER_US * 434;
		778: note_dur = CYCLES_PER_US * 103732;
		779: note_dur = CYCLES_PER_US * 434;
		780: note_dur = CYCLES_PER_US * 103732;
		781: note_dur = CYCLES_PER_US * 434;
		782: note_dur = CYCLES_PER_US * 103732;
		783: note_dur = CYCLES_PER_US * 434;
		784: note_dur = CYCLES_PER_US * 103732;
		785: note_dur = CYCLES_PER_US * 434;
		786: note_dur = CYCLES_PER_US * 103732;
		787: note_dur = CYCLES_PER_US * 434;
		788: note_dur = CYCLES_PER_US * 103732;
		789: note_dur = CYCLES_PER_US * 434;
		790: note_dur = CYCLES_PER_US * 103732;
		791: note_dur = CYCLES_PER_US * 434;
		792: note_dur = CYCLES_PER_US * 103732;
		793: note_dur = CYCLES_PER_US * 434;
		794: note_dur = CYCLES_PER_US * 103732;
		795: note_dur = CYCLES_PER_US * 434;
		796: note_dur = CYCLES_PER_US * 103732;
		797: note_dur = CYCLES_PER_US * 434;
		798: note_dur = CYCLES_PER_US * 103732;
		799: note_dur = CYCLES_PER_US * 434;
		800: note_dur = CYCLES_PER_US * 103732;
		801: note_dur = CYCLES_PER_US * 434;
		802: note_dur = CYCLES_PER_US * 103732;
		803: note_dur = CYCLES_PER_US * 434;
		804: note_dur = CYCLES_PER_US * 103732;
		805: note_dur = CYCLES_PER_US * 434;
		806: note_dur = CYCLES_PER_US * 103732;
		807: note_dur = CYCLES_PER_US * 434;
		808: note_dur = CYCLES_PER_US * 103732;
		809: note_dur = CYCLES_PER_US * 434;
		810: note_dur = CYCLES_PER_US * 103732;
		811: note_dur = CYCLES_PER_US * 434;
		812: note_dur = CYCLES_PER_US * 103732;
		813: note_dur = CYCLES_PER_US * 208767;
		814: note_dur = CYCLES_PER_US * 103732;
		815: note_dur = CYCLES_PER_US * 434;
		816: note_dur = CYCLES_PER_US * 103732;
		817: note_dur = CYCLES_PER_US * 434;
		818: note_dur = CYCLES_PER_US * 103732;
		819: note_dur = CYCLES_PER_US * 434;
		820: note_dur = CYCLES_PER_US * 103732;
		821: note_dur = CYCLES_PER_US * 434;
		822: note_dur = CYCLES_PER_US * 103732;
		823: note_dur = CYCLES_PER_US * 434;
		824: note_dur = CYCLES_PER_US * 103732;
		825: note_dur = CYCLES_PER_US * 434;
		826: note_dur = CYCLES_PER_US * 103732;
		827: note_dur = CYCLES_PER_US * 434;
		828: note_dur = CYCLES_PER_US * 103732;
		829: note_dur = CYCLES_PER_US * 434;
		830: note_dur = CYCLES_PER_US * 103732;
		831: note_dur = CYCLES_PER_US * 434;
		832: note_dur = CYCLES_PER_US * 103732;
		833: note_dur = CYCLES_PER_US * 434;
		834: note_dur = CYCLES_PER_US * 103732;
		835: note_dur = CYCLES_PER_US * 434;
		836: note_dur = CYCLES_PER_US * 103732;
		837: note_dur = CYCLES_PER_US * 434;
		838: note_dur = CYCLES_PER_US * 103732;
		839: note_dur = CYCLES_PER_US * 434;
		840: note_dur = CYCLES_PER_US * 103732;
		841: note_dur = CYCLES_PER_US * 434;
		842: note_dur = CYCLES_PER_US * 207899;
		843: note_dur = CYCLES_PER_US * 417100;
		844: note_dur = CYCLES_PER_US * 207899;
		845: note_dur = CYCLES_PER_US * 434;
		846: note_dur = CYCLES_PER_US * 103732;
		847: note_dur = CYCLES_PER_US * 434;
		848: note_dur = CYCLES_PER_US * 103732;
		849: note_dur = CYCLES_PER_US * 434;
		850: note_dur = CYCLES_PER_US * 103732;
		851: note_dur = CYCLES_PER_US * 434;
		852: note_dur = CYCLES_PER_US * 103732;
		853: note_dur = CYCLES_PER_US * 434;
		854: note_dur = CYCLES_PER_US * 103732;
		855: note_dur = CYCLES_PER_US * 434;
		856: note_dur = CYCLES_PER_US * 103732;
		857: note_dur = CYCLES_PER_US * 434;
		858: note_dur = CYCLES_PER_US * 103732;
		859: note_dur = CYCLES_PER_US * 434;
		860: note_dur = CYCLES_PER_US * 103732;
		861: note_dur = CYCLES_PER_US * 434;
		862: note_dur = CYCLES_PER_US * 103732;
		863: note_dur = CYCLES_PER_US * 434;
		864: note_dur = CYCLES_PER_US * 103732;
		865: note_dur = CYCLES_PER_US * 434;
		866: note_dur = CYCLES_PER_US * 103732;
		867: note_dur = CYCLES_PER_US * 434;
		868: note_dur = CYCLES_PER_US * 103732;
		869: note_dur = CYCLES_PER_US * 434;
		870: note_dur = CYCLES_PER_US * 103732;
		871: note_dur = CYCLES_PER_US * 434;
		872: note_dur = CYCLES_PER_US * 103732;
		873: note_dur = CYCLES_PER_US * 434;
		874: note_dur = CYCLES_PER_US * 103732;
		875: note_dur = CYCLES_PER_US * 434;
		876: note_dur = CYCLES_PER_US * 103732;
		877: note_dur = CYCLES_PER_US * 434;
		878: note_dur = CYCLES_PER_US * 103732;
		879: note_dur = CYCLES_PER_US * 434;
		880: note_dur = CYCLES_PER_US * 103732;
		881: note_dur = CYCLES_PER_US * 434;
		882: note_dur = CYCLES_PER_US * 103732;
		883: note_dur = CYCLES_PER_US * 434;
		884: note_dur = CYCLES_PER_US * 103732;
		885: note_dur = CYCLES_PER_US * 434;
		886: note_dur = CYCLES_PER_US * 103732;
		887: note_dur = CYCLES_PER_US * 434;
		888: note_dur = CYCLES_PER_US * 103732;
		889: note_dur = CYCLES_PER_US * 434;
		890: note_dur = CYCLES_PER_US * 103732;
		891: note_dur = CYCLES_PER_US * 434;
		892: note_dur = CYCLES_PER_US * 103732;
		893: note_dur = CYCLES_PER_US * 434;
		894: note_dur = CYCLES_PER_US * 103732;
		895: note_dur = CYCLES_PER_US * 434;
		896: note_dur = CYCLES_PER_US * 103732;
		897: note_dur = CYCLES_PER_US * 434;
		898: note_dur = CYCLES_PER_US * 312065;
		899: note_dur = CYCLES_PER_US * 434;
		900: note_dur = CYCLES_PER_US * 103732;
		901: note_dur = CYCLES_PER_US * 434;
		902: note_dur = CYCLES_PER_US * 207899;
		903: note_dur = CYCLES_PER_US * 434;
		904: note_dur = CYCLES_PER_US * 103732;
		905: note_dur = CYCLES_PER_US * 434;
		906: note_dur = CYCLES_PER_US * 51649;
		907: note_dur = CYCLES_PER_US * 434;
		908: note_dur = CYCLES_PER_US * 51649;
		909: note_dur = CYCLES_PER_US * 434;
		910: note_dur = CYCLES_PER_US * 207899;
		911: note_dur = CYCLES_PER_US * 312934;
		912: note_dur = CYCLES_PER_US * 103732;
		913: note_dur = CYCLES_PER_US * 434;
		914: note_dur = CYCLES_PER_US * 69010;
		915: note_dur = CYCLES_PER_US * 434;
		916: note_dur = CYCLES_PER_US * 69010;
		917: note_dur = CYCLES_PER_US * 434;
		918: note_dur = CYCLES_PER_US * 69010;
		919: note_dur = CYCLES_PER_US * 434;
		920: note_dur = CYCLES_PER_US * 207899;
		921: note_dur = CYCLES_PER_US * 434;
		922: note_dur = CYCLES_PER_US * 207899;
		923: note_dur = CYCLES_PER_US * 434;
		924: note_dur = CYCLES_PER_US * 312065;
		925: note_dur = CYCLES_PER_US * 434;
		926: note_dur = CYCLES_PER_US * 103732;
		927: note_dur = CYCLES_PER_US * 434;
		928: note_dur = CYCLES_PER_US * 103732;
		929: note_dur = CYCLES_PER_US * 434;
		930: note_dur = CYCLES_PER_US * 312065;
		931: note_dur = CYCLES_PER_US * 434;
		932: note_dur = CYCLES_PER_US * 0;
		933: note_dur = CYCLES_PER_US * 0;
		934: note_dur = CYCLES_PER_US * 0;
		935: note_dur = CYCLES_PER_US * 0;
		936: note_dur = CYCLES_PER_US * 416232;
		937: note_dur = CYCLES_PER_US * 0;
		938: note_dur = CYCLES_PER_US * 0;
		939: note_dur = CYCLES_PER_US * 0;
		940: note_dur = CYCLES_PER_US * 0;
		941: note_dur = CYCLES_PER_US * 434;
		942: note_dur = CYCLES_PER_US * 0;
		943: note_dur = CYCLES_PER_US * 0;
		944: note_dur = CYCLES_PER_US * 0;
		945: note_dur = CYCLES_PER_US * 103732;
		946: note_dur = CYCLES_PER_US * 0;
		947: note_dur = CYCLES_PER_US * 0;
		948: note_dur = CYCLES_PER_US * 0;
		949: note_dur = CYCLES_PER_US * 434;
		950: note_dur = CYCLES_PER_US * 103732;
		951: note_dur = CYCLES_PER_US * 434;
		952: note_dur = CYCLES_PER_US * 103732;
		953: note_dur = CYCLES_PER_US * 434;
		954: note_dur = CYCLES_PER_US * 103732;
		955: note_dur = CYCLES_PER_US * 434;
		956: note_dur = CYCLES_PER_US * 103732;
		957: note_dur = CYCLES_PER_US * 434;
		958: note_dur = CYCLES_PER_US * 103732;
		959: note_dur = CYCLES_PER_US * 434;
		960: note_dur = CYCLES_PER_US * 103732;
		961: note_dur = CYCLES_PER_US * 434;
		962: note_dur = CYCLES_PER_US * 103732;
		963: note_dur = CYCLES_PER_US * 434;
		964: note_dur = CYCLES_PER_US * 207899;
		965: note_dur = CYCLES_PER_US * 312934;
		966: note_dur = CYCLES_PER_US * 103732;
		967: note_dur = CYCLES_PER_US * 434;
		968: note_dur = CYCLES_PER_US * 103732;
		969: note_dur = CYCLES_PER_US * 434;
		970: note_dur = CYCLES_PER_US * 103732;
		971: note_dur = CYCLES_PER_US * 434;
		972: note_dur = CYCLES_PER_US * 312065;
		973: note_dur = CYCLES_PER_US * 434;
		974: note_dur = CYCLES_PER_US * 103732;
		975: note_dur = CYCLES_PER_US * 434;
		976: note_dur = CYCLES_PER_US * 0;
		977: note_dur = CYCLES_PER_US * 0;
		978: note_dur = CYCLES_PER_US * 0;
		979: note_dur = CYCLES_PER_US * 832898;
		980: note_dur = CYCLES_PER_US * 0;
		981: note_dur = CYCLES_PER_US * 0;
		982: note_dur = CYCLES_PER_US * 0;
		983: note_dur = CYCLES_PER_US * 434;
		984: note_dur = CYCLES_PER_US * 0;
		985: note_dur = CYCLES_PER_US * 0;
		986: note_dur = CYCLES_PER_US * 103732;
		987: note_dur = CYCLES_PER_US * 0;
		988: note_dur = CYCLES_PER_US * 0;
		989: note_dur = CYCLES_PER_US * 434;
		990: note_dur = CYCLES_PER_US * 103732;
		991: note_dur = CYCLES_PER_US * 434;
		992: note_dur = CYCLES_PER_US * 103732;
		993: note_dur = CYCLES_PER_US * 434;
		994: note_dur = CYCLES_PER_US * 103732;
		995: note_dur = CYCLES_PER_US * 434;
		996: note_dur = CYCLES_PER_US * 103732;
		997: note_dur = CYCLES_PER_US * 434;
		998: note_dur = CYCLES_PER_US * 103732;
		999: note_dur = CYCLES_PER_US * 434;
		1000: note_dur = CYCLES_PER_US * 103732;
		1001: note_dur = CYCLES_PER_US * 434;
		1002: note_dur = CYCLES_PER_US * 103732;
		1003: note_dur = CYCLES_PER_US * 434;
		1004: note_dur = CYCLES_PER_US * 103732;
		1005: note_dur = CYCLES_PER_US * 434;
		1006: note_dur = CYCLES_PER_US * 103732;
		1007: note_dur = CYCLES_PER_US * 434;
		1008: note_dur = CYCLES_PER_US * 103732;
		1009: note_dur = CYCLES_PER_US * 434;
		1010: note_dur = CYCLES_PER_US * 103732;
		1011: note_dur = CYCLES_PER_US * 434;
		1012: note_dur = CYCLES_PER_US * 103732;
		1013: note_dur = CYCLES_PER_US * 434;
		1014: note_dur = CYCLES_PER_US * 207899;
		1015: note_dur = CYCLES_PER_US * 434;
		1016: note_dur = CYCLES_PER_US * 103732;
		1017: note_dur = CYCLES_PER_US * 312934;
		1018: note_dur = CYCLES_PER_US * 51649;
		1019: note_dur = CYCLES_PER_US * 434;
		1020: note_dur = CYCLES_PER_US * 51649;
		1021: note_dur = CYCLES_PER_US * 434;
		1022: note_dur = CYCLES_PER_US * 207899;
		1023: note_dur = CYCLES_PER_US * 312934;
		1024: note_dur = CYCLES_PER_US * 103732;
		1025: note_dur = CYCLES_PER_US * 434;
		1026: note_dur = CYCLES_PER_US * 103732;
		1027: note_dur = CYCLES_PER_US * 434;
		1028: note_dur = CYCLES_PER_US * 103732;
		1029: note_dur = CYCLES_PER_US * 434;
		1030: note_dur = CYCLES_PER_US * 103732;
		1031: note_dur = CYCLES_PER_US * 434;
		1032: note_dur = CYCLES_PER_US * 103732;
		1033: note_dur = CYCLES_PER_US * 434;
		1034: note_dur = CYCLES_PER_US * 103732;
		1035: note_dur = CYCLES_PER_US * 434;
		1036: note_dur = CYCLES_PER_US * 103732;
		1037: note_dur = CYCLES_PER_US * 434;
		1038: note_dur = CYCLES_PER_US * 103732;
		1039: note_dur = CYCLES_PER_US * 434;
		1040: note_dur = CYCLES_PER_US * 103732;
		1041: note_dur = CYCLES_PER_US * 434;
		1042: note_dur = CYCLES_PER_US * 103732;
		1043: note_dur = CYCLES_PER_US * 434;
		1044: note_dur = CYCLES_PER_US * 103732;
		1045: note_dur = CYCLES_PER_US * 434;
		1046: note_dur = CYCLES_PER_US * 207899;
		1047: note_dur = CYCLES_PER_US * 434;
		1048: note_dur = CYCLES_PER_US * 103732;
		1049: note_dur = CYCLES_PER_US * 434;
		1050: note_dur = CYCLES_PER_US * 103732;
		1051: note_dur = CYCLES_PER_US * 434;
		1052: note_dur = CYCLES_PER_US * 103732;
		1053: note_dur = CYCLES_PER_US * 434;
		1054: note_dur = CYCLES_PER_US * 103732;
		1055: note_dur = CYCLES_PER_US * 434;
		1056: note_dur = CYCLES_PER_US * 103732;
		1057: note_dur = CYCLES_PER_US * 434;
		1058: note_dur = CYCLES_PER_US * 103732;
		1059: note_dur = CYCLES_PER_US * 434;
		1060: note_dur = CYCLES_PER_US * 103732;
		1061: note_dur = CYCLES_PER_US * 434;
		1062: note_dur = CYCLES_PER_US * 103732;
		1063: note_dur = CYCLES_PER_US * 434;
		1064: note_dur = CYCLES_PER_US * 103732;
		1065: note_dur = CYCLES_PER_US * 434;
		1066: note_dur = CYCLES_PER_US * 103732;
		1067: note_dur = CYCLES_PER_US * 434;
		1068: note_dur = CYCLES_PER_US * 103732;
		1069: note_dur = CYCLES_PER_US * 434;
		1070: note_dur = CYCLES_PER_US * 103732;
		1071: note_dur = CYCLES_PER_US * 434;
		1072: note_dur = CYCLES_PER_US * 103732;
		1073: note_dur = CYCLES_PER_US * 434;
		1074: note_dur = CYCLES_PER_US * 103732;
		1075: note_dur = CYCLES_PER_US * 434;
		1076: note_dur = CYCLES_PER_US * 103732;
		1077: note_dur = CYCLES_PER_US * 434;
		1078: note_dur = CYCLES_PER_US * 103732;
		1079: note_dur = CYCLES_PER_US * 434;
		1080: note_dur = CYCLES_PER_US * 103732;
		1081: note_dur = CYCLES_PER_US * 434;
		1082: note_dur = CYCLES_PER_US * 103732;
		1083: note_dur = CYCLES_PER_US * 434;
		1084: note_dur = CYCLES_PER_US * 103732;
		1085: note_dur = CYCLES_PER_US * 434;
		1086: note_dur = CYCLES_PER_US * 103732;
		1087: note_dur = CYCLES_PER_US * 434;
		1088: note_dur = CYCLES_PER_US * 103732;
		1089: note_dur = CYCLES_PER_US * 434;
		1090: note_dur = CYCLES_PER_US * 103732;
		1091: note_dur = CYCLES_PER_US * 434;
		1092: note_dur = CYCLES_PER_US * 103732;
		1093: note_dur = CYCLES_PER_US * 434;
		1094: note_dur = CYCLES_PER_US * 103732;
		1095: note_dur = CYCLES_PER_US * 434;
		1096: note_dur = CYCLES_PER_US * 103732;
		1097: note_dur = CYCLES_PER_US * 434;
		1098: note_dur = CYCLES_PER_US * 103732;
		1099: note_dur = CYCLES_PER_US * 104601;
		1100: note_dur = CYCLES_PER_US * 0;
		1101: note_dur = CYCLES_PER_US * 103732;
		1102: note_dur = CYCLES_PER_US * 0;
		1103: note_dur = CYCLES_PER_US * 434;
		1104: note_dur = CYCLES_PER_US * 69010;
		1105: note_dur = CYCLES_PER_US * 434;
		1106: note_dur = CYCLES_PER_US * 69010;
		1107: note_dur = CYCLES_PER_US * 434;
		1108: note_dur = CYCLES_PER_US * 69010;
		1109: note_dur = CYCLES_PER_US * 434;
		1110: note_dur = CYCLES_PER_US * 207899;
		1111: note_dur = CYCLES_PER_US * 434;
		1112: note_dur = CYCLES_PER_US * 103732;
		1113: note_dur = CYCLES_PER_US * 434;
		1114: note_dur = CYCLES_PER_US * 416232;
		1115: note_dur = CYCLES_PER_US * 434;
		1116: note_dur = CYCLES_PER_US * 103732;
		1117: note_dur = CYCLES_PER_US * 434;
		1118: note_dur = CYCLES_PER_US * 103732;
		1119: note_dur = CYCLES_PER_US * 434;
		1120: note_dur = CYCLES_PER_US * 103732;
		1121: note_dur = CYCLES_PER_US * 312934;
		1122: note_dur = CYCLES_PER_US * 103732;
		1123: note_dur = CYCLES_PER_US * 434;
		1124: note_dur = CYCLES_PER_US * 69010;
		1125: note_dur = CYCLES_PER_US * 434;
		1126: note_dur = CYCLES_PER_US * 69010;
		1127: note_dur = CYCLES_PER_US * 434;
		1128: note_dur = CYCLES_PER_US * 69010;
		1129: note_dur = CYCLES_PER_US * 434;
		1130: note_dur = CYCLES_PER_US * 103732;
		1131: note_dur = CYCLES_PER_US * 434;
		1132: note_dur = CYCLES_PER_US * 520398;
		1133: note_dur = CYCLES_PER_US * 520398;
		default: note_dur = 0;
	endcase
end
endmodule