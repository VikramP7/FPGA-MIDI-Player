module song4_pitch(
	input logic [10:0] note_index,
	output logic [6:0] note_pitch
);

always_comb begin
	case (note_index)
		0: note_pitch = 66;
		1: note_pitch = 0;
		2: note_pitch = 62;
		3: note_pitch = 0;
		4: note_pitch = 59;
		5: note_pitch = 0;
		6: note_pitch = 55;
		7: note_pitch = 0;
		8: note_pitch = 58;
		9: note_pitch = 0;
		10: note_pitch = 59;
		11: note_pitch = 0;
		12: note_pitch = 57;
		13: note_pitch = 0;
		14: note_pitch = 62;
		15: note_pitch = 0;
		16: note_pitch = 58;
		17: note_pitch = 0;
		18: note_pitch = 55;
		19: note_pitch = 0;
		20: note_pitch = 51;
		21: note_pitch = 0;
		22: note_pitch = 54;
		23: note_pitch = 0;
		24: note_pitch = 55;
		25: note_pitch = 0;
		26: note_pitch = 53;
		27: note_pitch = 0;
		28: note_pitch = 58;
		29: note_pitch = 0;
		30: note_pitch = 59;
		31: note_pitch = 0;
		32: note_pitch = 57;
		33: note_pitch = 0;
		34: note_pitch = 62;
		35: note_pitch = 0;
		36: note_pitch = 63;
		37: note_pitch = 0;
		38: note_pitch = 63;
		39: note_pitch = 0;
		40: note_pitch = 66;
		41: note_pitch = 0;
		42: note_pitch = 67;
		43: note_pitch = 0;
		44: note_pitch = 67;
		45: note_pitch = 0;
		46: note_pitch = 70;
		47: note_pitch = 0;
		48: note_pitch = 66;
		49: note_pitch = 0;
		50: note_pitch = 66;
		51: note_pitch = 0;
		52: note_pitch = 66;
		53: note_pitch = 0;
		54: note_pitch = 62;
		55: note_pitch = 0;
		56: note_pitch = 59;
		57: note_pitch = 0;
		58: note_pitch = 55;
		59: note_pitch = 0;
		60: note_pitch = 58;
		61: note_pitch = 0;
		62: note_pitch = 59;
		63: note_pitch = 0;
		64: note_pitch = 57;
		65: note_pitch = 0;
		66: note_pitch = 62;
		67: note_pitch = 0;
		68: note_pitch = 58;
		69: note_pitch = 0;
		70: note_pitch = 55;
		71: note_pitch = 0;
		72: note_pitch = 51;
		73: note_pitch = 0;
		74: note_pitch = 54;
		75: note_pitch = 0;
		76: note_pitch = 55;
		77: note_pitch = 0;
		78: note_pitch = 53;
		79: note_pitch = 0;
		80: note_pitch = 58;
		81: note_pitch = 0;
		82: note_pitch = 59;
		83: note_pitch = 0;
		84: note_pitch = 57;
		85: note_pitch = 0;
		86: note_pitch = 62;
		87: note_pitch = 0;
		88: note_pitch = 63;
		89: note_pitch = 0;
		90: note_pitch = 63;
		91: note_pitch = 0;
		92: note_pitch = 66;
		93: note_pitch = 0;
		94: note_pitch = 67;
		95: note_pitch = 0;
		96: note_pitch = 67;
		97: note_pitch = 0;
		98: note_pitch = 70;
		99: note_pitch = 0;
		100: note_pitch = 61;
		101: note_pitch = 0;
		102: note_pitch = 64;
		103: note_pitch = 0;
		104: note_pitch = 68;
		105: note_pitch = 0;
		106: note_pitch = 71;
		107: note_pitch = 0;
		108: note_pitch = 70;
		109: note_pitch = 0;
		110: note_pitch = 68;
		111: note_pitch = 0;
		112: note_pitch = 66;
		113: note_pitch = 0;
		114: note_pitch = 63;
		115: note_pitch = 0;
		116: note_pitch = 59;
		117: note_pitch = 0;
		118: note_pitch = 62;
		119: note_pitch = 0;
		120: note_pitch = 64;
		121: note_pitch = 0;
		122: note_pitch = 66;
		123: note_pitch = 0;
		124: note_pitch = 69;
		125: note_pitch = 0;
		126: note_pitch = 67;
		127: note_pitch = 0;
		128: note_pitch = 62;
		129: note_pitch = 0;
		130: note_pitch = 59;
		131: note_pitch = 0;
		132: note_pitch = 60;
		133: note_pitch = 0;
		134: note_pitch = 56;
		135: note_pitch = 0;
		136: note_pitch = 55;
		137: note_pitch = 0;
		138: note_pitch = 53;
		139: note_pitch = 0;
		140: note_pitch = 51;
		141: note_pitch = 0;
		142: note_pitch = 53;
		143: note_pitch = 0;
		144: note_pitch = 55;
		145: note_pitch = 0;
		146: note_pitch = 56;
		147: note_pitch = 0;
		148: note_pitch = 58;
		149: note_pitch = 0;
		150: note_pitch = 60;
		151: note_pitch = 0;
		152: note_pitch = 62;
		153: note_pitch = 0;
		154: note_pitch = 63;
		155: note_pitch = 0;
		156: note_pitch = 64;
		157: note_pitch = 0;
		158: note_pitch = 60;
		159: note_pitch = 0;
		160: note_pitch = 57;
		161: note_pitch = 0;
		162: note_pitch = 55;
		163: note_pitch = 0;
		164: note_pitch = 54;
		165: note_pitch = 0;
		166: note_pitch = 63;
		167: note_pitch = 0;
		168: note_pitch = 62;
		169: note_pitch = 0;
		170: note_pitch = 60;
		171: note_pitch = 0;
		172: note_pitch = 59;
		173: note_pitch = 0;
		174: note_pitch = 62;
		175: note_pitch = 0;
		176: note_pitch = 67;
		177: note_pitch = 0;
		178: note_pitch = 71;
		179: note_pitch = 0;
		180: note_pitch = 62;
		181: note_pitch = 0;
		182: note_pitch = 65;
		183: note_pitch = 0;
		184: note_pitch = 68;
		185: note_pitch = 0;
		186: note_pitch = 72;
		187: note_pitch = 0;
		188: note_pitch = 63;
		189: note_pitch = 0;
		190: note_pitch = 65;
		191: note_pitch = 0;
		192: note_pitch = 67;
		193: note_pitch = 0;
		194: note_pitch = 70;
		195: note_pitch = 0;
		196: note_pitch = 64;
		197: note_pitch = 0;
		198: note_pitch = 68;
		199: note_pitch = 0;
		200: note_pitch = 70;
		201: note_pitch = 0;
		202: note_pitch = 73;
		203: note_pitch = 0;
		204: note_pitch = 70;
		205: note_pitch = 0;
		206: note_pitch = 68;
		207: note_pitch = 0;
		208: note_pitch = 66;
		209: note_pitch = 0;
		210: note_pitch = 70;
		211: note_pitch = 0;
		212: note_pitch = 69;
		213: note_pitch = 0;
		214: note_pitch = 68;
		215: note_pitch = 0;
		216: note_pitch = 67;
		217: note_pitch = 0;
		218: note_pitch = 65;
		219: note_pitch = 0;
		220: note_pitch = 63;
		221: note_pitch = 0;
		222: note_pitch = 62;
		223: note_pitch = 0;
		224: note_pitch = 60;
		225: note_pitch = 0;
		226: note_pitch = 58;
		227: note_pitch = 0;
		228: note_pitch = 68;
		229: note_pitch = 0;
		230: note_pitch = 67;
		231: note_pitch = 0;
		232: note_pitch = 62;
		233: note_pitch = 0;
		234: note_pitch = 65;
		235: note_pitch = 0;
		236: note_pitch = 63;
		237: note_pitch = 0;
		238: note_pitch = 62;
		239: note_pitch = 0;
		240: note_pitch = 65;
		241: note_pitch = 0;
		242: note_pitch = 64;
		243: note_pitch = 0;
		244: note_pitch = 60;
		245: note_pitch = 0;
		246: note_pitch = 57;
		247: note_pitch = 0;
		248: note_pitch = 52;
		249: note_pitch = 0;
		250: note_pitch = 55;
		251: note_pitch = 0;
		252: note_pitch = 52;
		253: note_pitch = 0;
		254: note_pitch = 54;
		255: note_pitch = 0;
		256: note_pitch = 63;
		257: note_pitch = 0;
		258: note_pitch = 62;
		259: note_pitch = 0;
		260: note_pitch = 60;
		261: note_pitch = 0;
		262: note_pitch = 59;
		263: note_pitch = 0;
		264: note_pitch = 57;
		265: note_pitch = 0;
		266: note_pitch = 55;
		267: note_pitch = 0;
		268: note_pitch = 57;
		269: note_pitch = 0;
		270: note_pitch = 59;
		271: note_pitch = 0;
		272: note_pitch = 62;
		273: note_pitch = 0;
		274: note_pitch = 63;
		275: note_pitch = 0;
		276: note_pitch = 61;
		277: note_pitch = 0;
		278: note_pitch = 59;
		279: note_pitch = 0;
		280: note_pitch = 58;
		281: note_pitch = 0;
		282: note_pitch = 54;
		283: note_pitch = 0;
		284: note_pitch = 56;
		285: note_pitch = 0;
		286: note_pitch = 58;
		287: note_pitch = 0;
		288: note_pitch = 59;
		289: note_pitch = 0;
		290: note_pitch = 61;
		291: note_pitch = 0;
		292: note_pitch = 63;
		293: note_pitch = 0;
		294: note_pitch = 66;
		295: note_pitch = 0;
		296: note_pitch = 70;
		297: note_pitch = 0;
		298: note_pitch = 69;
		299: note_pitch = 0;
		300: note_pitch = 68;
		301: note_pitch = 0;
		302: note_pitch = 67;
		303: note_pitch = 0;
		304: note_pitch = 65;
		305: note_pitch = 0;
		306: note_pitch = 67;
		307: note_pitch = 0;
		308: note_pitch = 66;
		309: note_pitch = 0;
		310: note_pitch = 65;
		311: note_pitch = 0;
		312: note_pitch = 62;
		313: note_pitch = 0;
		314: note_pitch = 63;
		315: note_pitch = 0;
		316: note_pitch = 65;
		317: note_pitch = 0;
		318: note_pitch = 67;
		319: note_pitch = 0;
		320: note_pitch = 70;
		321: note_pitch = 0;
		322: note_pitch = 75;
		323: note_pitch = 0;
		324: note_pitch = 70;
		325: note_pitch = 0;
		326: note_pitch = 70;
		327: note_pitch = 0;
		328: note_pitch = 71;
		329: note_pitch = 0;
		330: note_pitch = 70;
		331: note_pitch = 0;
		332: note_pitch = 66;
		333: note_pitch = 0;
		334: note_pitch = 71;
		335: note_pitch = 72;
		336: note_pitch = 73;
		337: note_pitch = 74;
		338: note_pitch = 0;
		339: note_pitch = 0;
		340: note_pitch = 0;
		341: note_pitch = 0;
		342: note_pitch = 72;
		343: note_pitch = 0;
		344: note_pitch = 71;
		345: note_pitch = 0;
		346: note_pitch = 62;
		347: note_pitch = 0;
		348: note_pitch = 67;
		349: note_pitch = 0;
		350: note_pitch = 71;
		351: note_pitch = 0;
		352: note_pitch = 70;
		353: note_pitch = 0;
		354: note_pitch = 69;
		355: note_pitch = 0;
		356: note_pitch = 68;
		357: note_pitch = 0;
		358: note_pitch = 72;
		359: note_pitch = 0;
		360: note_pitch = 70;
		361: note_pitch = 0;
		362: note_pitch = 67;
		363: note_pitch = 0;
		364: note_pitch = 65;
		365: note_pitch = 0;
		366: note_pitch = 63;
		367: note_pitch = 0;
		368: note_pitch = 67;
		369: note_pitch = 0;
		370: note_pitch = 63;
		371: note_pitch = 0;
		372: note_pitch = 70;
		373: note_pitch = 71;
		374: note_pitch = 72;
		375: note_pitch = 73;
		376: note_pitch = 74;
		377: note_pitch = 0;
		378: note_pitch = 0;
		379: note_pitch = 0;
		380: note_pitch = 0;
		381: note_pitch = 0;
		382: note_pitch = 70;
		383: note_pitch = 0;
		384: note_pitch = 66;
		385: note_pitch = 0;
		386: note_pitch = 62;
		387: note_pitch = 0;
		388: note_pitch = 62;
		389: note_pitch = 0;
		390: note_pitch = 67;
		391: note_pitch = 0;
		392: note_pitch = 71;
		393: note_pitch = 0;
		394: note_pitch = 62;
		395: note_pitch = 0;
		396: note_pitch = 65;
		397: note_pitch = 0;
		398: note_pitch = 68;
		399: note_pitch = 0;
		400: note_pitch = 72;
		401: note_pitch = 0;
		402: note_pitch = 63;
		403: note_pitch = 0;
		404: note_pitch = 65;
		405: note_pitch = 0;
		406: note_pitch = 67;
		407: note_pitch = 0;
		408: note_pitch = 70;
		409: note_pitch = 0;
		410: note_pitch = 64;
		411: note_pitch = 0;
		412: note_pitch = 66;
		413: note_pitch = 0;
		414: note_pitch = 68;
		415: note_pitch = 0;
		416: note_pitch = 70;
		417: note_pitch = 0;
		418: note_pitch = 66;
		419: note_pitch = 0;
		420: note_pitch = 63;
		421: note_pitch = 0;
		422: note_pitch = 61;
		423: note_pitch = 0;
		424: note_pitch = 59;
		425: note_pitch = 0;
		426: note_pitch = 58;
		427: note_pitch = 0;
		428: note_pitch = 54;
		429: note_pitch = 0;
		430: note_pitch = 60;
		431: note_pitch = 0;
		432: note_pitch = 62;
		433: note_pitch = 0;
		434: note_pitch = 63;
		435: note_pitch = 0;
		436: note_pitch = 60;
		437: note_pitch = 0;
		438: note_pitch = 67;
		439: note_pitch = 0;
		440: note_pitch = 65;
		441: note_pitch = 0;
		442: note_pitch = 62;
		443: note_pitch = 0;
		444: note_pitch = 60;
		445: note_pitch = 0;
		446: note_pitch = 58;
		447: note_pitch = 0;
		448: note_pitch = 68;
		449: note_pitch = 0;
		450: note_pitch = 67;
		451: note_pitch = 0;
		452: note_pitch = 63;
		453: note_pitch = 0;
		454: note_pitch = 57;
		455: note_pitch = 0;
		456: note_pitch = 60;
		457: note_pitch = 0;
		458: note_pitch = 64;
		459: note_pitch = 0;
		460: note_pitch = 71;
		461: note_pitch = 0;
		462: note_pitch = 69;
		463: note_pitch = 0;
		464: note_pitch = 66;
		465: note_pitch = 0;
		466: note_pitch = 64;
		467: note_pitch = 0;
		468: note_pitch = 62;
		469: note_pitch = 0;
		470: note_pitch = 64;
		471: note_pitch = 0;
		472: note_pitch = 66;
		473: note_pitch = 0;
		474: note_pitch = 69;
		475: note_pitch = 0;
		476: note_pitch = 67;
		477: note_pitch = 0;
		478: note_pitch = 69;
		479: note_pitch = 0;
		480: note_pitch = 71;
		481: note_pitch = 0;
		482: note_pitch = 70;
		483: note_pitch = 0;
		484: note_pitch = 71;
		485: note_pitch = 0;
		486: note_pitch = 70;
		487: note_pitch = 0;
		488: note_pitch = 66;
		489: note_pitch = 0;
		490: note_pitch = 68;
		491: note_pitch = 0;
		492: note_pitch = 70;
		493: note_pitch = 0;
		494: note_pitch = 66;
		495: note_pitch = 0;
		496: note_pitch = 63;
		497: note_pitch = 0;
		498: note_pitch = 61;
		499: note_pitch = 0;
		500: note_pitch = 59;
		501: note_pitch = 0;
		502: note_pitch = 60;
		503: note_pitch = 0;
		504: note_pitch = 62;
		505: note_pitch = 0;
		506: note_pitch = 63;
		507: note_pitch = 0;
		508: note_pitch = 60;
		509: note_pitch = 0;
		510: note_pitch = 67;
		511: note_pitch = 0;
		512: note_pitch = 65;
		513: note_pitch = 0;
		514: note_pitch = 62;
		515: note_pitch = 0;
		516: note_pitch = 58;
		517: note_pitch = 0;
		518: note_pitch = 58;
		519: note_pitch = 0;
		520: note_pitch = 67;
		521: note_pitch = 0;
		522: note_pitch = 61;
		523: note_pitch = 0;
		524: note_pitch = 64;
		525: note_pitch = 0;
		526: note_pitch = 68;
		527: note_pitch = 0;
		528: note_pitch = 71;
		529: note_pitch = 0;
		530: note_pitch = 66;
		531: note_pitch = 0;
		532: note_pitch = 68;
		533: note_pitch = 0;
		534: note_pitch = 70;
		535: note_pitch = 0;
		536: note_pitch = 73;
		537: note_pitch = 0;
		538: note_pitch = 59;
		539: note_pitch = 66;
		540: note_pitch = 0;
		541: note_pitch = 0;
		542: note_pitch = 61;
		543: note_pitch = 0;
		544: note_pitch = 63;
		545: note_pitch = 0;
		546: note_pitch = 66;
		547: note_pitch = 0;
		548: note_pitch = 62;
		549: note_pitch = 0;
		550: note_pitch = 64;
		551: note_pitch = 0;
		552: note_pitch = 66;
		553: note_pitch = 0;
		554: note_pitch = 69;
		555: note_pitch = 0;
		556: note_pitch = 67;
		557: note_pitch = 0;
		558: note_pitch = 62;
		559: note_pitch = 0;
		560: note_pitch = 59;
		561: note_pitch = 0;
		562: note_pitch = 60;
		563: note_pitch = 0;
		564: note_pitch = 56;
		565: note_pitch = 0;
		566: note_pitch = 55;
		567: note_pitch = 0;
		568: note_pitch = 53;
		569: note_pitch = 0;
		570: note_pitch = 51;
		571: note_pitch = 0;
		572: note_pitch = 53;
		573: note_pitch = 0;
		574: note_pitch = 55;
		575: note_pitch = 0;
		576: note_pitch = 56;
		577: note_pitch = 0;
		578: note_pitch = 58;
		579: note_pitch = 0;
		580: note_pitch = 60;
		581: note_pitch = 0;
		582: note_pitch = 62;
		583: note_pitch = 0;
		584: note_pitch = 65;
		585: note_pitch = 0;
		586: note_pitch = 64;
		587: note_pitch = 0;
		588: note_pitch = 68;
		589: note_pitch = 0;
		590: note_pitch = 71;
		591: note_pitch = 0;
		592: note_pitch = 62;
		593: note_pitch = 0;
		594: note_pitch = 64;
		595: note_pitch = 0;
		596: note_pitch = 66;
		597: note_pitch = 0;
		598: note_pitch = 67;
		599: note_pitch = 0;
		600: note_pitch = 69;
		601: note_pitch = 0;
		602: note_pitch = 71;
		603: note_pitch = 0;
		604: note_pitch = 74;
		605: note_pitch = 0;
		606: note_pitch = 68;
		607: note_pitch = 0;
		608: note_pitch = 72;
		609: note_pitch = 0;
		610: note_pitch = 70;
		611: note_pitch = 0;
		612: note_pitch = 68;
		613: note_pitch = 0;
		614: note_pitch = 67;
		615: note_pitch = 0;
		616: note_pitch = 63;
		617: note_pitch = 0;
		618: note_pitch = 65;
		619: note_pitch = 0;
		620: note_pitch = 67;
		621: note_pitch = 0;
		622: note_pitch = 64;
		623: note_pitch = 0;
		624: note_pitch = 66;
		625: note_pitch = 0;
		626: note_pitch = 68;
		627: note_pitch = 0;
		628: note_pitch = 70;
		629: note_pitch = 0;
		630: note_pitch = 73;
		631: note_pitch = 0;
		632: note_pitch = 70;
		633: note_pitch = 0;
		634: note_pitch = 68;
		635: note_pitch = 0;
		636: note_pitch = 66;
		637: note_pitch = 0;
		638: note_pitch = 63;
		639: note_pitch = 0;
		640: note_pitch = 70;
		641: note_pitch = 71;
		642: note_pitch = 72;
		643: note_pitch = 73;
		644: note_pitch = 74;
		645: note_pitch = 0;
		646: note_pitch = 0;
		647: note_pitch = 0;
		648: note_pitch = 0;
		649: note_pitch = 0;
		650: note_pitch = 72;
		651: note_pitch = 0;
		652: note_pitch = 71;
		653: note_pitch = 0;
		654: note_pitch = 70;
		655: note_pitch = 0;
		656: note_pitch = 68;
		657: note_pitch = 0;
		658: note_pitch = 67;
		659: note_pitch = 0;
		660: note_pitch = 65;
		661: note_pitch = 0;
		662: note_pitch = 63;
		663: note_pitch = 0;
		664: note_pitch = 65;
		665: note_pitch = 0;
		666: note_pitch = 67;
		667: note_pitch = 0;
		668: note_pitch = 70;
		669: note_pitch = 0;
		670: note_pitch = 71;
		671: note_pitch = 72;
		672: note_pitch = 73;
		673: note_pitch = 74;
		674: note_pitch = 0;
		675: note_pitch = 0;
		676: note_pitch = 0;
		677: note_pitch = 0;
		678: note_pitch = 74;
		679: note_pitch = 0;
		680: note_pitch = 73;
		681: note_pitch = 0;
		682: note_pitch = 74;
		683: note_pitch = 0;
		684: note_pitch = 71;
		685: note_pitch = 0;
		686: note_pitch = 67;
		687: note_pitch = 0;
		688: note_pitch = 69;
		689: note_pitch = 0;
		690: note_pitch = 66;
		691: note_pitch = 0;
		692: note_pitch = 67;
		693: note_pitch = 0;
		694: note_pitch = 62;
		695: note_pitch = 0;
		696: note_pitch = 59;
		697: note_pitch = 0;
		698: note_pitch = 55;
		699: note_pitch = 0;
		700: note_pitch = 63;
		701: note_pitch = 0;
		702: note_pitch = 59;
		703: note_pitch = 0;
		704: note_pitch = 58;
		705: note_pitch = 0;
		706: note_pitch = 54;
		707: note_pitch = 0;
		708: note_pitch = 56;
		709: note_pitch = 0;
		710: note_pitch = 54;
		711: note_pitch = 0;
		712: note_pitch = 56;
		713: note_pitch = 0;
		714: note_pitch = 58;
		715: note_pitch = 0;
		716: note_pitch = 59;
		717: note_pitch = 0;
		718: note_pitch = 61;
		719: note_pitch = 0;
		720: note_pitch = 63;
		721: note_pitch = 0;
		722: note_pitch = 66;
		723: note_pitch = 0;
		724: note_pitch = 70;
		725: note_pitch = 0;
		726: note_pitch = 66;
		727: note_pitch = 0;
		728: note_pitch = 63;
		729: note_pitch = 0;
		730: note_pitch = 59;
		731: note_pitch = 0;
		732: note_pitch = 68;
		733: note_pitch = 0;
		734: note_pitch = 67;
		735: note_pitch = 0;
		736: note_pitch = 66;
		737: note_pitch = 0;
		738: note_pitch = 65;
		739: note_pitch = 0;
		740: note_pitch = 63;
		741: note_pitch = 0;
		742: note_pitch = 62;
		743: note_pitch = 0;
		744: note_pitch = 60;
		745: note_pitch = 0;
		746: note_pitch = 58;
		747: note_pitch = 0;
		748: note_pitch = 56;
		749: note_pitch = 0;
		750: note_pitch = 55;
		751: note_pitch = 0;
		752: note_pitch = 53;
		753: note_pitch = 0;
		754: note_pitch = 51;
		755: note_pitch = 0;
		756: note_pitch = 53;
		757: note_pitch = 0;
		758: note_pitch = 55;
		759: note_pitch = 0;
		760: note_pitch = 58;
		761: note_pitch = 0;
		762: note_pitch = 63;
		763: note_pitch = 0;
		764: note_pitch = 54;
		765: note_pitch = 0;
		766: note_pitch = 59;
		767: note_pitch = 0;
		768: note_pitch = 63;
		769: note_pitch = 0;
		770: note_pitch = 62;
		771: note_pitch = 0;
		772: note_pitch = 64;
		773: note_pitch = 0;
		774: note_pitch = 66;
		775: note_pitch = 0;
		776: note_pitch = 69;
		777: note_pitch = 0;
		778: note_pitch = 67;
		779: note_pitch = 0;
		780: note_pitch = 62;
		781: note_pitch = 0;
		782: note_pitch = 59;
		783: note_pitch = 0;
		784: note_pitch = 55;
		785: note_pitch = 0;
		786: note_pitch = 60;
		787: note_pitch = 0;
		788: note_pitch = 56;
		789: note_pitch = 0;
		790: note_pitch = 55;
		791: note_pitch = 0;
		792: note_pitch = 53;
		793: note_pitch = 0;
		794: note_pitch = 51;
		795: note_pitch = 0;
		796: note_pitch = 53;
		797: note_pitch = 0;
		798: note_pitch = 55;
		799: note_pitch = 0;
		800: note_pitch = 56;
		801: note_pitch = 0;
		802: note_pitch = 58;
		803: note_pitch = 0;
		804: note_pitch = 60;
		805: note_pitch = 0;
		806: note_pitch = 62;
		807: note_pitch = 0;
		808: note_pitch = 65;
		809: note_pitch = 0;
		810: note_pitch = 64;
		811: note_pitch = 0;
		812: note_pitch = 68;
		813: note_pitch = 0;
		814: note_pitch = 71;
		815: note_pitch = 0;
		816: note_pitch = 62;
		817: note_pitch = 0;
		818: note_pitch = 64;
		819: note_pitch = 0;
		820: note_pitch = 69;
		821: note_pitch = 0;
		822: note_pitch = 67;
		823: note_pitch = 0;
		824: note_pitch = 69;
		825: note_pitch = 0;
		826: note_pitch = 71;
		827: note_pitch = 0;
		828: note_pitch = 72;
		829: note_pitch = 0;
		830: note_pitch = 62;
		831: note_pitch = 0;
		832: note_pitch = 65;
		833: note_pitch = 0;
		834: note_pitch = 68;
		835: note_pitch = 0;
		836: note_pitch = 72;
		837: note_pitch = 0;
		838: note_pitch = 63;
		839: note_pitch = 0;
		840: note_pitch = 65;
		841: note_pitch = 0;
		842: note_pitch = 67;
		843: note_pitch = 0;
		844: note_pitch = 66;
		845: note_pitch = 0;
		846: note_pitch = 63;
		847: note_pitch = 0;
		848: note_pitch = 61;
		849: note_pitch = 0;
		850: note_pitch = 59;
		851: note_pitch = 0;
		852: note_pitch = 61;
		853: note_pitch = 0;
		854: note_pitch = 63;
		855: note_pitch = 0;
		856: note_pitch = 66;
		857: note_pitch = 0;
		858: note_pitch = 70;
		859: note_pitch = 0;
		860: note_pitch = 69;
		861: note_pitch = 0;
		862: note_pitch = 68;
		863: note_pitch = 0;
		864: note_pitch = 67;
		865: note_pitch = 0;
		866: note_pitch = 65;
		867: note_pitch = 0;
		868: note_pitch = 63;
		869: note_pitch = 0;
		870: note_pitch = 62;
		871: note_pitch = 0;
		872: note_pitch = 60;
		873: note_pitch = 0;
		874: note_pitch = 60;
		875: note_pitch = 0;
		876: note_pitch = 68;
		877: note_pitch = 0;
		878: note_pitch = 67;
		879: note_pitch = 0;
		880: note_pitch = 62;
		881: note_pitch = 0;
		882: note_pitch = 65;
		883: note_pitch = 0;
		884: note_pitch = 63;
		885: note_pitch = 0;
		886: note_pitch = 60;
		887: note_pitch = 0;
		888: note_pitch = 65;
		889: note_pitch = 0;
		890: note_pitch = 64;
		891: note_pitch = 0;
		892: note_pitch = 60;
		893: note_pitch = 0;
		894: note_pitch = 57;
		895: note_pitch = 0;
		896: note_pitch = 52;
		897: note_pitch = 0;
		898: note_pitch = 55;
		899: note_pitch = 0;
		900: note_pitch = 54;
		901: note_pitch = 0;
		902: note_pitch = 62;
		903: note_pitch = 0;
		904: note_pitch = 59;
		905: note_pitch = 0;
		906: note_pitch = 62;
		907: note_pitch = 0;
		908: note_pitch = 67;
		909: note_pitch = 0;
		910: note_pitch = 71;
		911: note_pitch = 0;
		912: note_pitch = 61;
		913: note_pitch = 0;
		914: note_pitch = 64;
		915: note_pitch = 0;
		916: note_pitch = 68;
		917: note_pitch = 0;
		918: note_pitch = 71;
		919: note_pitch = 0;
		920: note_pitch = 70;
		921: note_pitch = 0;
		922: note_pitch = 73;
		923: note_pitch = 0;
		924: note_pitch = 73;
		925: note_pitch = 0;
		926: note_pitch = 70;
		927: note_pitch = 0;
		928: note_pitch = 66;
		929: note_pitch = 0;
		930: note_pitch = 63;
		931: note_pitch = 0;
		932: note_pitch = 70;
		933: note_pitch = 71;
		934: note_pitch = 72;
		935: note_pitch = 73;
		936: note_pitch = 74;
		937: note_pitch = 0;
		938: note_pitch = 0;
		939: note_pitch = 0;
		940: note_pitch = 0;
		941: note_pitch = 0;
		942: note_pitch = 73;
		943: note_pitch = 72;
		944: note_pitch = 71;
		945: note_pitch = 70;
		946: note_pitch = 0;
		947: note_pitch = 0;
		948: note_pitch = 0;
		949: note_pitch = 0;
		950: note_pitch = 68;
		951: note_pitch = 0;
		952: note_pitch = 67;
		953: note_pitch = 0;
		954: note_pitch = 63;
		955: note_pitch = 0;
		956: note_pitch = 63;
		957: note_pitch = 0;
		958: note_pitch = 65;
		959: note_pitch = 0;
		960: note_pitch = 67;
		961: note_pitch = 0;
		962: note_pitch = 70;
		963: note_pitch = 0;
		964: note_pitch = 75;
		965: note_pitch = 0;
		966: note_pitch = 75;
		967: note_pitch = 0;
		968: note_pitch = 73;
		969: note_pitch = 0;
		970: note_pitch = 71;
		971: note_pitch = 0;
		972: note_pitch = 70;
		973: note_pitch = 0;
		974: note_pitch = 66;
		975: note_pitch = 0;
		976: note_pitch = 71;
		977: note_pitch = 72;
		978: note_pitch = 73;
		979: note_pitch = 74;
		980: note_pitch = 0;
		981: note_pitch = 0;
		982: note_pitch = 0;
		983: note_pitch = 0;
		984: note_pitch = 73;
		985: note_pitch = 72;
		986: note_pitch = 71;
		987: note_pitch = 0;
		988: note_pitch = 0;
		989: note_pitch = 0;
		990: note_pitch = 62;
		991: note_pitch = 0;
		992: note_pitch = 67;
		993: note_pitch = 0;
		994: note_pitch = 71;
		995: note_pitch = 0;
		996: note_pitch = 70;
		997: note_pitch = 0;
		998: note_pitch = 69;
		999: note_pitch = 0;
		1000: note_pitch = 68;
		1001: note_pitch = 0;
		1002: note_pitch = 72;
		1003: note_pitch = 0;
		1004: note_pitch = 70;
		1005: note_pitch = 0;
		1006: note_pitch = 67;
		1007: note_pitch = 0;
		1008: note_pitch = 65;
		1009: note_pitch = 0;
		1010: note_pitch = 63;
		1011: note_pitch = 0;
		1012: note_pitch = 67;
		1013: note_pitch = 0;
		1014: note_pitch = 70;
		1015: note_pitch = 0;
		1016: note_pitch = 75;
		1017: note_pitch = 0;
		1018: note_pitch = 67;
		1019: note_pitch = 0;
		1020: note_pitch = 71;
		1021: note_pitch = 0;
		1022: note_pitch = 69;
		1023: note_pitch = 0;
		1024: note_pitch = 62;
		1025: note_pitch = 0;
		1026: note_pitch = 67;
		1027: note_pitch = 0;
		1028: note_pitch = 71;
		1029: note_pitch = 0;
		1030: note_pitch = 62;
		1031: note_pitch = 0;
		1032: note_pitch = 63;
		1033: note_pitch = 0;
		1034: note_pitch = 68;
		1035: note_pitch = 0;
		1036: note_pitch = 72;
		1037: note_pitch = 0;
		1038: note_pitch = 63;
		1039: note_pitch = 0;
		1040: note_pitch = 65;
		1041: note_pitch = 0;
		1042: note_pitch = 67;
		1043: note_pitch = 0;
		1044: note_pitch = 70;
		1045: note_pitch = 0;
		1046: note_pitch = 75;
		1047: note_pitch = 0;
		1048: note_pitch = 73;
		1049: note_pitch = 0;
		1050: note_pitch = 71;
		1051: note_pitch = 0;
		1052: note_pitch = 70;
		1053: note_pitch = 0;
		1054: note_pitch = 68;
		1055: note_pitch = 0;
		1056: note_pitch = 66;
		1057: note_pitch = 0;
		1058: note_pitch = 64;
		1059: note_pitch = 0;
		1060: note_pitch = 63;
		1061: note_pitch = 0;
		1062: note_pitch = 61;
		1063: note_pitch = 0;
		1064: note_pitch = 59;
		1065: note_pitch = 0;
		1066: note_pitch = 54;
		1067: note_pitch = 0;
		1068: note_pitch = 60;
		1069: note_pitch = 0;
		1070: note_pitch = 62;
		1071: note_pitch = 0;
		1072: note_pitch = 63;
		1073: note_pitch = 0;
		1074: note_pitch = 65;
		1075: note_pitch = 0;
		1076: note_pitch = 67;
		1077: note_pitch = 0;
		1078: note_pitch = 65;
		1079: note_pitch = 0;
		1080: note_pitch = 62;
		1081: note_pitch = 0;
		1082: note_pitch = 60;
		1083: note_pitch = 0;
		1084: note_pitch = 58;
		1085: note_pitch = 0;
		1086: note_pitch = 68;
		1087: note_pitch = 0;
		1088: note_pitch = 67;
		1089: note_pitch = 0;
		1090: note_pitch = 62;
		1091: note_pitch = 0;
		1092: note_pitch = 65;
		1093: note_pitch = 0;
		1094: note_pitch = 63;
		1095: note_pitch = 0;
		1096: note_pitch = 62;
		1097: note_pitch = 0;
		1098: note_pitch = 60;
		1099: note_pitch = 0;
		1100: note_pitch = 57;
		1101: note_pitch = 64;
		1102: note_pitch = 0;
		1103: note_pitch = 0;
		1104: note_pitch = 60;
		1105: note_pitch = 0;
		1106: note_pitch = 64;
		1107: note_pitch = 0;
		1108: note_pitch = 67;
		1109: note_pitch = 0;
		1110: note_pitch = 71;
		1111: note_pitch = 0;
		1112: note_pitch = 67;
		1113: note_pitch = 0;
		1114: note_pitch = 71;
		1115: note_pitch = 0;
		1116: note_pitch = 67;
		1117: note_pitch = 0;
		1118: note_pitch = 71;
		1119: note_pitch = 0;
		1120: note_pitch = 74;
		1121: note_pitch = 0;
		1122: note_pitch = 61;
		1123: note_pitch = 0;
		1124: note_pitch = 64;
		1125: note_pitch = 0;
		1126: note_pitch = 68;
		1127: note_pitch = 0;
		1128: note_pitch = 71;
		1129: note_pitch = 0;
		1130: note_pitch = 70;
		1131: note_pitch = 0;
		1132: note_pitch = 73;
		1133: note_pitch = 0;
		default: note_pitch = 0;
	endcase
end
endmodule