module song5_pitch(
	input logic [10:0] note_index,
	output logic [6:0] note_pitch
);

always_comb begin
	case (note_index)
		0: note_pitch = 58;
		1: note_pitch = 0;
		2: note_pitch = 63;
		3: note_pitch = 0;
		4: note_pitch = 66;
		5: note_pitch = 0;
		6: note_pitch = 68;
		7: note_pitch = 0;
		8: note_pitch = 69;
		9: note_pitch = 0;
		10: note_pitch = 70;
		11: note_pitch = 0;
		12: note_pitch = 69;
		13: note_pitch = 0;
		14: note_pitch = 68;
		15: note_pitch = 0;
		16: note_pitch = 66;
		17: note_pitch = 0;
		18: note_pitch = 58;
		19: note_pitch = 0;
		20: note_pitch = 59;
		21: note_pitch = 0;
		22: note_pitch = 60;
		23: note_pitch = 0;
		24: note_pitch = 61;
		25: note_pitch = 0;
		26: note_pitch = 63;
		27: note_pitch = 0;
		28: note_pitch = 65;
		29: note_pitch = 0;
		30: note_pitch = 66;
		31: note_pitch = 0;
		32: note_pitch = 65;
		33: note_pitch = 0;
		34: note_pitch = 63;
		35: note_pitch = 0;
		36: note_pitch = 61;
		37: note_pitch = 0;
		38: note_pitch = 63;
		39: note_pitch = 0;
		40: note_pitch = 61;
		41: note_pitch = 0;
		42: note_pitch = 63;
		43: note_pitch = 0;
		44: note_pitch = 61;
		45: note_pitch = 0;
		46: note_pitch = 58;
		47: note_pitch = 0;
		48: note_pitch = 56;
		49: note_pitch = 0;
		50: note_pitch = 58;
		51: note_pitch = 0;
		52: note_pitch = 58;
		53: note_pitch = 0;
		54: note_pitch = 63;
		55: note_pitch = 0;
		56: note_pitch = 66;
		57: note_pitch = 0;
		58: note_pitch = 68;
		59: note_pitch = 0;
		60: note_pitch = 69;
		61: note_pitch = 0;
		62: note_pitch = 70;
		63: note_pitch = 0;
		64: note_pitch = 69;
		65: note_pitch = 0;
		66: note_pitch = 68;
		67: note_pitch = 0;
		68: note_pitch = 66;
		69: note_pitch = 0;
		70: note_pitch = 58;
		71: note_pitch = 0;
		72: note_pitch = 59;
		73: note_pitch = 0;
		74: note_pitch = 60;
		75: note_pitch = 0;
		76: note_pitch = 61;
		77: note_pitch = 0;
		78: note_pitch = 63;
		79: note_pitch = 0;
		80: note_pitch = 61;
		81: note_pitch = 0;
		82: note_pitch = 63;
		83: note_pitch = 0;
		84: note_pitch = 61;
		85: note_pitch = 0;
		86: note_pitch = 58;
		87: note_pitch = 0;
		88: note_pitch = 56;
		89: note_pitch = 0;
		90: note_pitch = 58;
		91: note_pitch = 0;
		92: note_pitch = 65;
		93: note_pitch = 0;
		94: note_pitch = 66;
		95: note_pitch = 0;
		96: note_pitch = 65;
		97: note_pitch = 0;
		98: note_pitch = 63;
		99: note_pitch = 0;
		100: note_pitch = 61;
		101: note_pitch = 0;
		102: note_pitch = 63;
		103: note_pitch = 0;
		104: note_pitch = 75;
		105: note_pitch = 0;
		106: note_pitch = 78;
		107: note_pitch = 0;
		108: note_pitch = 75;
		109: note_pitch = 0;
		110: note_pitch = 71;
		111: note_pitch = 0;
		112: note_pitch = 68;
		113: note_pitch = 0;
		114: note_pitch = 70;
		115: note_pitch = 0;
		116: note_pitch = 71;
		117: note_pitch = 0;
		118: note_pitch = 72;
		119: note_pitch = 0;
		120: note_pitch = 73;
		121: note_pitch = 0;
		122: note_pitch = 77;
		123: note_pitch = 0;
		124: note_pitch = 73;
		125: note_pitch = 0;
		126: note_pitch = 70;
		127: note_pitch = 0;
		128: note_pitch = 66;
		129: note_pitch = 0;
		130: note_pitch = 68;
		131: note_pitch = 0;
		132: note_pitch = 69;
		133: note_pitch = 0;
		134: note_pitch = 70;
		135: note_pitch = 0;
		136: note_pitch = 71;
		137: note_pitch = 0;
		138: note_pitch = 75;
		139: note_pitch = 0;
		140: note_pitch = 71;
		141: note_pitch = 0;
		142: note_pitch = 68;
		143: note_pitch = 0;
		144: note_pitch = 65;
		145: note_pitch = 0;
		146: note_pitch = 66;
		147: note_pitch = 0;
		148: note_pitch = 68;
		149: note_pitch = 0;
		150: note_pitch = 69;
		151: note_pitch = 0;
		152: note_pitch = 70;
		153: note_pitch = 0;
		154: note_pitch = 69;
		155: note_pitch = 0;
		156: note_pitch = 70;
		157: note_pitch = 0;
		158: note_pitch = 71;
		159: note_pitch = 0;
		160: note_pitch = 73;
		161: note_pitch = 0;
		162: note_pitch = 73;
		163: note_pitch = 0;
		164: note_pitch = 72;
		165: note_pitch = 0;
		166: note_pitch = 73;
		167: note_pitch = 0;
		168: note_pitch = 74;
		169: note_pitch = 0;
		170: note_pitch = 75;
		171: note_pitch = 0;
		172: note_pitch = 78;
		173: note_pitch = 0;
		174: note_pitch = 75;
		175: note_pitch = 0;
		176: note_pitch = 71;
		177: note_pitch = 0;
		178: note_pitch = 68;
		179: note_pitch = 0;
		180: note_pitch = 70;
		181: note_pitch = 0;
		182: note_pitch = 72;
		183: note_pitch = 0;
		184: note_pitch = 73;
		185: note_pitch = 0;
		186: note_pitch = 77;
		187: note_pitch = 0;
		188: note_pitch = 73;
		189: note_pitch = 0;
		190: note_pitch = 70;
		191: note_pitch = 0;
		192: note_pitch = 66;
		193: note_pitch = 0;
		194: note_pitch = 68;
		195: note_pitch = 0;
		196: note_pitch = 69;
		197: note_pitch = 0;
		198: note_pitch = 70;
		199: note_pitch = 0;
		200: note_pitch = 71;
		201: note_pitch = 0;
		202: note_pitch = 75;
		203: note_pitch = 0;
		204: note_pitch = 71;
		205: note_pitch = 0;
		206: note_pitch = 68;
		207: note_pitch = 0;
		208: note_pitch = 65;
		209: note_pitch = 0;
		210: note_pitch = 68;
		211: note_pitch = 0;
		212: note_pitch = 73;
		213: note_pitch = 0;
		214: note_pitch = 71;
		215: note_pitch = 0;
		216: note_pitch = 70;
		217: note_pitch = 0;
		218: note_pitch = 58;
		219: note_pitch = 0;
		220: note_pitch = 63;
		221: note_pitch = 0;
		222: note_pitch = 66;
		223: note_pitch = 0;
		224: note_pitch = 68;
		225: note_pitch = 0;
		226: note_pitch = 69;
		227: note_pitch = 0;
		228: note_pitch = 70;
		229: note_pitch = 0;
		230: note_pitch = 69;
		231: note_pitch = 0;
		232: note_pitch = 68;
		233: note_pitch = 0;
		234: note_pitch = 66;
		235: note_pitch = 0;
		236: note_pitch = 58;
		237: note_pitch = 0;
		238: note_pitch = 59;
		239: note_pitch = 0;
		240: note_pitch = 60;
		241: note_pitch = 0;
		242: note_pitch = 61;
		243: note_pitch = 0;
		244: note_pitch = 63;
		245: note_pitch = 0;
		246: note_pitch = 65;
		247: note_pitch = 0;
		248: note_pitch = 66;
		249: note_pitch = 0;
		250: note_pitch = 65;
		251: note_pitch = 0;
		252: note_pitch = 63;
		253: note_pitch = 0;
		254: note_pitch = 61;
		255: note_pitch = 0;
		256: note_pitch = 63;
		257: note_pitch = 0;
		258: note_pitch = 61;
		259: note_pitch = 0;
		260: note_pitch = 63;
		261: note_pitch = 0;
		262: note_pitch = 61;
		263: note_pitch = 0;
		264: note_pitch = 58;
		265: note_pitch = 0;
		266: note_pitch = 56;
		267: note_pitch = 0;
		268: note_pitch = 58;
		269: note_pitch = 0;
		270: note_pitch = 58;
		271: note_pitch = 0;
		272: note_pitch = 63;
		273: note_pitch = 0;
		274: note_pitch = 66;
		275: note_pitch = 0;
		276: note_pitch = 68;
		277: note_pitch = 0;
		278: note_pitch = 69;
		279: note_pitch = 0;
		280: note_pitch = 70;
		281: note_pitch = 0;
		282: note_pitch = 69;
		283: note_pitch = 0;
		284: note_pitch = 68;
		285: note_pitch = 0;
		286: note_pitch = 66;
		287: note_pitch = 0;
		288: note_pitch = 58;
		289: note_pitch = 0;
		290: note_pitch = 59;
		291: note_pitch = 0;
		292: note_pitch = 60;
		293: note_pitch = 0;
		294: note_pitch = 61;
		295: note_pitch = 0;
		296: note_pitch = 63;
		297: note_pitch = 0;
		298: note_pitch = 65;
		299: note_pitch = 0;
		300: note_pitch = 66;
		301: note_pitch = 0;
		302: note_pitch = 65;
		303: note_pitch = 0;
		304: note_pitch = 63;
		305: note_pitch = 0;
		306: note_pitch = 61;
		307: note_pitch = 0;
		308: note_pitch = 63;
		309: note_pitch = 0;
		310: note_pitch = 61;
		311: note_pitch = 0;
		312: note_pitch = 63;
		313: note_pitch = 0;
		314: note_pitch = 61;
		315: note_pitch = 0;
		316: note_pitch = 58;
		317: note_pitch = 0;
		318: note_pitch = 56;
		319: note_pitch = 0;
		320: note_pitch = 58;
		321: note_pitch = 0;
		322: note_pitch = 68;
		323: note_pitch = 70;
		324: note_pitch = 0;
		325: note_pitch = 0;
		326: note_pitch = 63;
		327: note_pitch = 0;
		328: note_pitch = 60;
		329: note_pitch = 0;
		330: note_pitch = 58;
		331: note_pitch = 0;
		332: note_pitch = 63;
		333: note_pitch = 0;
		334: note_pitch = 65;
		335: note_pitch = 0;
		336: note_pitch = 66;
		337: note_pitch = 0;
		338: note_pitch = 75;
		339: note_pitch = 0;
		340: note_pitch = 70;
		341: note_pitch = 0;
		342: note_pitch = 68;
		343: note_pitch = 0;
		344: note_pitch = 66;
		345: note_pitch = 0;
		346: note_pitch = 68;
		347: note_pitch = 0;
		348: note_pitch = 63;
		349: note_pitch = 0;
		350: note_pitch = 66;
		351: note_pitch = 0;
		352: note_pitch = 63;
		353: note_pitch = 0;
		354: note_pitch = 65;
		355: note_pitch = 0;
		356: note_pitch = 66;
		357: note_pitch = 0;
		358: note_pitch = 70;
		359: note_pitch = 0;
		360: note_pitch = 63;
		361: note_pitch = 0;
		362: note_pitch = 66;
		363: note_pitch = 0;
		364: note_pitch = 63;
		365: note_pitch = 0;
		366: note_pitch = 65;
		367: note_pitch = 0;
		368: note_pitch = 68;
		369: note_pitch = 0;
		370: note_pitch = 63;
		371: note_pitch = 0;
		372: note_pitch = 66;
		373: note_pitch = 0;
		374: note_pitch = 63;
		375: note_pitch = 0;
		376: note_pitch = 65;
		377: note_pitch = 0;
		378: note_pitch = 61;
		379: note_pitch = 0;
		380: note_pitch = 58;
		381: note_pitch = 0;
		382: note_pitch = 56;
		383: note_pitch = 0;
		384: note_pitch = 63;
		385: note_pitch = 0;
		386: note_pitch = 66;
		387: note_pitch = 0;
		388: note_pitch = 63;
		389: note_pitch = 0;
		390: note_pitch = 65;
		391: note_pitch = 0;
		392: note_pitch = 68;
		393: note_pitch = 0;
		394: note_pitch = 63;
		395: note_pitch = 0;
		396: note_pitch = 66;
		397: note_pitch = 0;
		398: note_pitch = 63;
		399: note_pitch = 0;
		400: note_pitch = 65;
		401: note_pitch = 0;
		402: note_pitch = 70;
		403: note_pitch = 0;
		404: note_pitch = 68;
		405: note_pitch = 0;
		406: note_pitch = 66;
		407: note_pitch = 0;
		408: note_pitch = 65;
		409: note_pitch = 0;
		410: note_pitch = 63;
		411: note_pitch = 0;
		412: note_pitch = 56;
		413: note_pitch = 0;
		414: note_pitch = 68;
		415: note_pitch = 0;
		416: note_pitch = 73;
		417: note_pitch = 0;
		418: note_pitch = 70;
		419: note_pitch = 0;
		420: note_pitch = 66;
		421: note_pitch = 0;
		422: note_pitch = 63;
		423: note_pitch = 0;
		424: note_pitch = 56;
		425: note_pitch = 0;
		426: note_pitch = 63;
		427: note_pitch = 0;
		428: note_pitch = 65;
		429: note_pitch = 0;
		430: note_pitch = 63;
		431: note_pitch = 0;
		432: note_pitch = 68;
		433: note_pitch = 0;
		434: note_pitch = 63;
		435: note_pitch = 0;
		436: note_pitch = 65;
		437: note_pitch = 0;
		438: note_pitch = 61;
		439: note_pitch = 0;
		440: note_pitch = 63;
		441: note_pitch = 0;
		442: note_pitch = 65;
		443: note_pitch = 0;
		444: note_pitch = 66;
		445: note_pitch = 0;
		446: note_pitch = 68;
		447: note_pitch = 0;
		448: note_pitch = 70;
		449: note_pitch = 0;
		450: note_pitch = 72;
		451: note_pitch = 0;
		452: note_pitch = 68;
		453: note_pitch = 0;
		454: note_pitch = 70;
		455: note_pitch = 0;
		456: note_pitch = 75;
		457: note_pitch = 0;
		458: note_pitch = 70;
		459: note_pitch = 0;
		460: note_pitch = 72;
		461: note_pitch = 0;
		462: note_pitch = 68;
		463: note_pitch = 0;
		464: note_pitch = 70;
		465: note_pitch = 0;
		466: note_pitch = 72;
		467: note_pitch = 0;
		468: note_pitch = 73;
		469: note_pitch = 0;
		470: note_pitch = 75;
		471: note_pitch = 76;
		472: note_pitch = 0;
		473: note_pitch = 77;
		474: note_pitch = 0;
		475: note_pitch = 76;
		476: note_pitch = 0;
		477: note_pitch = 77;
		478: note_pitch = 0;
		479: note_pitch = 0;
		480: note_pitch = 73;
		481: note_pitch = 0;
		482: note_pitch = 70;
		483: note_pitch = 0;
		484: note_pitch = 66;
		485: note_pitch = 0;
		486: note_pitch = 75;
		487: note_pitch = 0;
		488: note_pitch = 71;
		489: note_pitch = 0;
		490: note_pitch = 68;
		491: note_pitch = 0;
		492: note_pitch = 73;
		493: note_pitch = 0;
		494: note_pitch = 70;
		495: note_pitch = 0;
		496: note_pitch = 66;
		497: note_pitch = 0;
		498: note_pitch = 65;
		499: note_pitch = 0;
		500: note_pitch = 61;
		501: note_pitch = 0;
		502: note_pitch = 63;
		503: note_pitch = 0;
		504: note_pitch = 65;
		505: note_pitch = 0;
		506: note_pitch = 66;
		507: note_pitch = 0;
		508: note_pitch = 68;
		509: note_pitch = 0;
		510: note_pitch = 70;
		511: note_pitch = 0;
		512: note_pitch = 63;
		513: note_pitch = 0;
		514: note_pitch = 63;
		515: note_pitch = 0;
		516: note_pitch = 56;
		517: note_pitch = 0;
		518: note_pitch = 68;
		519: note_pitch = 0;
		520: note_pitch = 56;
		521: note_pitch = 0;
		522: note_pitch = 66;
		523: note_pitch = 0;
		524: note_pitch = 65;
		525: note_pitch = 0;
		526: note_pitch = 63;
		527: note_pitch = 0;
		528: note_pitch = 56;
		529: note_pitch = 0;
		530: note_pitch = 68;
		531: note_pitch = 0;
		532: note_pitch = 63;
		533: note_pitch = 0;
		534: note_pitch = 65;
		535: note_pitch = 0;
		536: note_pitch = 66;
		537: note_pitch = 0;
		538: note_pitch = 56;
		539: note_pitch = 0;
		540: note_pitch = 68;
		541: note_pitch = 0;
		542: note_pitch = 63;
		543: note_pitch = 0;
		544: note_pitch = 66;
		545: note_pitch = 0;
		546: note_pitch = 65;
		547: note_pitch = 0;
		548: note_pitch = 63;
		549: note_pitch = 0;
		550: note_pitch = 56;
		551: note_pitch = 0;
		552: note_pitch = 65;
		553: note_pitch = 0;
		554: note_pitch = 61;
		555: note_pitch = 0;
		556: note_pitch = 63;
		557: note_pitch = 0;
		558: note_pitch = 59;
		559: note_pitch = 0;
		560: note_pitch = 58;
		561: note_pitch = 0;
		562: note_pitch = 58;
		563: note_pitch = 0;
		564: note_pitch = 63;
		565: note_pitch = 0;
		566: note_pitch = 66;
		567: note_pitch = 0;
		568: note_pitch = 68;
		569: note_pitch = 0;
		570: note_pitch = 58;
		571: note_pitch = 0;
		572: note_pitch = 58;
		573: note_pitch = 0;
		574: note_pitch = 63;
		575: note_pitch = 0;
		576: note_pitch = 66;
		577: note_pitch = 0;
		578: note_pitch = 68;
		579: note_pitch = 0;
		580: note_pitch = 69;
		581: note_pitch = 0;
		582: note_pitch = 70;
		583: note_pitch = 0;
		584: note_pitch = 69;
		585: note_pitch = 0;
		586: note_pitch = 68;
		587: note_pitch = 0;
		588: note_pitch = 66;
		589: note_pitch = 0;
		590: note_pitch = 58;
		591: note_pitch = 0;
		592: note_pitch = 59;
		593: note_pitch = 0;
		594: note_pitch = 60;
		595: note_pitch = 0;
		596: note_pitch = 61;
		597: note_pitch = 0;
		598: note_pitch = 63;
		599: note_pitch = 0;
		600: note_pitch = 65;
		601: note_pitch = 0;
		602: note_pitch = 66;
		603: note_pitch = 0;
		604: note_pitch = 65;
		605: note_pitch = 0;
		606: note_pitch = 63;
		607: note_pitch = 0;
		608: note_pitch = 61;
		609: note_pitch = 0;
		610: note_pitch = 63;
		611: note_pitch = 0;
		612: note_pitch = 61;
		613: note_pitch = 0;
		614: note_pitch = 63;
		615: note_pitch = 0;
		616: note_pitch = 61;
		617: note_pitch = 0;
		618: note_pitch = 58;
		619: note_pitch = 0;
		620: note_pitch = 56;
		621: note_pitch = 0;
		622: note_pitch = 58;
		623: note_pitch = 0;
		624: note_pitch = 58;
		625: note_pitch = 0;
		626: note_pitch = 63;
		627: note_pitch = 0;
		628: note_pitch = 66;
		629: note_pitch = 0;
		630: note_pitch = 68;
		631: note_pitch = 0;
		632: note_pitch = 69;
		633: note_pitch = 0;
		634: note_pitch = 70;
		635: note_pitch = 0;
		636: note_pitch = 69;
		637: note_pitch = 0;
		638: note_pitch = 68;
		639: note_pitch = 0;
		640: note_pitch = 66;
		641: note_pitch = 0;
		642: note_pitch = 58;
		643: note_pitch = 0;
		644: note_pitch = 59;
		645: note_pitch = 0;
		646: note_pitch = 60;
		647: note_pitch = 0;
		648: note_pitch = 61;
		649: note_pitch = 0;
		650: note_pitch = 63;
		651: note_pitch = 0;
		652: note_pitch = 61;
		653: note_pitch = 0;
		654: note_pitch = 63;
		655: note_pitch = 0;
		656: note_pitch = 61;
		657: note_pitch = 0;
		658: note_pitch = 58;
		659: note_pitch = 0;
		660: note_pitch = 56;
		661: note_pitch = 0;
		662: note_pitch = 58;
		663: note_pitch = 0;
		664: note_pitch = 65;
		665: note_pitch = 0;
		666: note_pitch = 66;
		667: note_pitch = 0;
		668: note_pitch = 65;
		669: note_pitch = 0;
		670: note_pitch = 63;
		671: note_pitch = 0;
		672: note_pitch = 61;
		673: note_pitch = 0;
		674: note_pitch = 63;
		675: note_pitch = 0;
		676: note_pitch = 75;
		677: note_pitch = 0;
		678: note_pitch = 78;
		679: note_pitch = 0;
		680: note_pitch = 75;
		681: note_pitch = 0;
		682: note_pitch = 71;
		683: note_pitch = 0;
		684: note_pitch = 68;
		685: note_pitch = 0;
		686: note_pitch = 70;
		687: note_pitch = 0;
		688: note_pitch = 71;
		689: note_pitch = 0;
		690: note_pitch = 72;
		691: note_pitch = 0;
		692: note_pitch = 73;
		693: note_pitch = 0;
		694: note_pitch = 77;
		695: note_pitch = 0;
		696: note_pitch = 73;
		697: note_pitch = 0;
		698: note_pitch = 70;
		699: note_pitch = 0;
		700: note_pitch = 66;
		701: note_pitch = 0;
		702: note_pitch = 68;
		703: note_pitch = 0;
		704: note_pitch = 69;
		705: note_pitch = 0;
		706: note_pitch = 70;
		707: note_pitch = 0;
		708: note_pitch = 71;
		709: note_pitch = 0;
		710: note_pitch = 75;
		711: note_pitch = 0;
		712: note_pitch = 71;
		713: note_pitch = 0;
		714: note_pitch = 68;
		715: note_pitch = 0;
		716: note_pitch = 65;
		717: note_pitch = 0;
		718: note_pitch = 66;
		719: note_pitch = 0;
		720: note_pitch = 68;
		721: note_pitch = 0;
		722: note_pitch = 69;
		723: note_pitch = 0;
		724: note_pitch = 70;
		725: note_pitch = 0;
		726: note_pitch = 69;
		727: note_pitch = 0;
		728: note_pitch = 70;
		729: note_pitch = 0;
		730: note_pitch = 71;
		731: note_pitch = 0;
		732: note_pitch = 73;
		733: note_pitch = 0;
		734: note_pitch = 73;
		735: note_pitch = 0;
		736: note_pitch = 72;
		737: note_pitch = 0;
		738: note_pitch = 73;
		739: note_pitch = 0;
		740: note_pitch = 74;
		741: note_pitch = 0;
		742: note_pitch = 75;
		743: note_pitch = 0;
		744: note_pitch = 78;
		745: note_pitch = 0;
		746: note_pitch = 75;
		747: note_pitch = 0;
		748: note_pitch = 71;
		749: note_pitch = 0;
		750: note_pitch = 68;
		751: note_pitch = 0;
		752: note_pitch = 70;
		753: note_pitch = 0;
		754: note_pitch = 72;
		755: note_pitch = 0;
		756: note_pitch = 73;
		757: note_pitch = 0;
		758: note_pitch = 77;
		759: note_pitch = 0;
		760: note_pitch = 73;
		761: note_pitch = 0;
		762: note_pitch = 70;
		763: note_pitch = 0;
		764: note_pitch = 66;
		765: note_pitch = 0;
		766: note_pitch = 68;
		767: note_pitch = 0;
		768: note_pitch = 69;
		769: note_pitch = 0;
		770: note_pitch = 70;
		771: note_pitch = 0;
		772: note_pitch = 71;
		773: note_pitch = 0;
		774: note_pitch = 75;
		775: note_pitch = 0;
		776: note_pitch = 71;
		777: note_pitch = 0;
		778: note_pitch = 68;
		779: note_pitch = 0;
		780: note_pitch = 65;
		781: note_pitch = 0;
		782: note_pitch = 68;
		783: note_pitch = 0;
		784: note_pitch = 73;
		785: note_pitch = 0;
		786: note_pitch = 71;
		787: note_pitch = 0;
		788: note_pitch = 70;
		789: note_pitch = 0;
		790: note_pitch = 58;
		791: note_pitch = 0;
		792: note_pitch = 63;
		793: note_pitch = 0;
		794: note_pitch = 66;
		795: note_pitch = 0;
		796: note_pitch = 68;
		797: note_pitch = 0;
		798: note_pitch = 69;
		799: note_pitch = 0;
		800: note_pitch = 70;
		801: note_pitch = 0;
		802: note_pitch = 69;
		803: note_pitch = 0;
		804: note_pitch = 68;
		805: note_pitch = 0;
		806: note_pitch = 66;
		807: note_pitch = 0;
		808: note_pitch = 58;
		809: note_pitch = 0;
		810: note_pitch = 59;
		811: note_pitch = 0;
		812: note_pitch = 60;
		813: note_pitch = 0;
		814: note_pitch = 61;
		815: note_pitch = 0;
		816: note_pitch = 63;
		817: note_pitch = 0;
		818: note_pitch = 65;
		819: note_pitch = 0;
		820: note_pitch = 66;
		821: note_pitch = 0;
		822: note_pitch = 65;
		823: note_pitch = 0;
		824: note_pitch = 63;
		825: note_pitch = 0;
		826: note_pitch = 61;
		827: note_pitch = 0;
		828: note_pitch = 63;
		829: note_pitch = 0;
		830: note_pitch = 61;
		831: note_pitch = 0;
		832: note_pitch = 63;
		833: note_pitch = 0;
		834: note_pitch = 61;
		835: note_pitch = 0;
		836: note_pitch = 58;
		837: note_pitch = 0;
		838: note_pitch = 56;
		839: note_pitch = 0;
		840: note_pitch = 58;
		841: note_pitch = 0;
		842: note_pitch = 58;
		843: note_pitch = 0;
		844: note_pitch = 63;
		845: note_pitch = 0;
		846: note_pitch = 66;
		847: note_pitch = 0;
		848: note_pitch = 68;
		849: note_pitch = 0;
		850: note_pitch = 69;
		851: note_pitch = 0;
		852: note_pitch = 70;
		853: note_pitch = 0;
		854: note_pitch = 69;
		855: note_pitch = 0;
		856: note_pitch = 68;
		857: note_pitch = 0;
		858: note_pitch = 66;
		859: note_pitch = 0;
		860: note_pitch = 58;
		861: note_pitch = 0;
		862: note_pitch = 59;
		863: note_pitch = 0;
		864: note_pitch = 60;
		865: note_pitch = 0;
		866: note_pitch = 61;
		867: note_pitch = 0;
		868: note_pitch = 63;
		869: note_pitch = 0;
		870: note_pitch = 61;
		871: note_pitch = 0;
		872: note_pitch = 63;
		873: note_pitch = 0;
		874: note_pitch = 61;
		875: note_pitch = 0;
		876: note_pitch = 58;
		877: note_pitch = 0;
		878: note_pitch = 56;
		879: note_pitch = 0;
		880: note_pitch = 58;
		881: note_pitch = 0;
		882: note_pitch = 65;
		883: note_pitch = 0;
		884: note_pitch = 66;
		885: note_pitch = 0;
		886: note_pitch = 65;
		887: note_pitch = 0;
		888: note_pitch = 63;
		889: note_pitch = 0;
		890: note_pitch = 61;
		891: note_pitch = 0;
		892: note_pitch = 63;
		893: note_pitch = 0;
		894: note_pitch = 61;
		895: note_pitch = 0;
		896: note_pitch = 63;
		897: note_pitch = 0;
		898: note_pitch = 61;
		899: note_pitch = 0;
		900: note_pitch = 58;
		901: note_pitch = 0;
		902: note_pitch = 56;
		903: note_pitch = 0;
		904: note_pitch = 58;
		905: note_pitch = 0;
		906: note_pitch = 61;
		907: note_pitch = 0;
		908: note_pitch = 63;
		909: note_pitch = 0;
		910: note_pitch = 61;
		911: note_pitch = 0;
		912: note_pitch = 58;
		913: note_pitch = 0;
		914: note_pitch = 56;
		915: note_pitch = 0;
		916: note_pitch = 58;
		917: note_pitch = 0;
		918: note_pitch = 65;
		919: note_pitch = 0;
		920: note_pitch = 66;
		921: note_pitch = 0;
		922: note_pitch = 65;
		923: note_pitch = 0;
		924: note_pitch = 63;
		925: note_pitch = 0;
		926: note_pitch = 61;
		927: note_pitch = 0;
		928: note_pitch = 63;
		929: note_pitch = 0;
		default: note_pitch = 0;
	endcase
end
endmodule