module song6_dur #(
	parameter int CLOCK_FREQ = 100_000_000
) (
	input logic [10:0] note_index,
	output logic [28:0] note_dur // max 10s at 100MHz clock
);

localparam real TEMPO_BPM = 120;
localparam real CYCLES_PER_BEAT = CLOCK_FREQ*(60/TEMPO_BPM);
localparam real CYCLES_PER_US = CLOCK_FREQ/1000_000;

always_comb begin
	// the quarter note is one beat and therfore can be multipled by CYCLES_PER_BEAT
	case (note_index)
		0: note_dur = CYCLES_PER_US * 170714;
		1: note_dur = CYCLES_PER_US * 714;
		2: note_dur = CYCLES_PER_US * 342143;
		3: note_dur = CYCLES_PER_US * 714;
		4: note_dur = CYCLES_PER_US * 170714;
		5: note_dur = CYCLES_PER_US * 714;
		6: note_dur = CYCLES_PER_US * 170714;
		7: note_dur = CYCLES_PER_US * 714;
		8: note_dur = CYCLES_PER_US * 170714;
		9: note_dur = CYCLES_PER_US * 172143;
		10: note_dur = CYCLES_PER_US * 170714;
		11: note_dur = CYCLES_PER_US * 714;
		12: note_dur = CYCLES_PER_US * 170714;
		13: note_dur = CYCLES_PER_US * 172143;
		14: note_dur = CYCLES_PER_US * 170714;
		15: note_dur = CYCLES_PER_US * 857857;
		16: note_dur = CYCLES_PER_US * 170714;
		17: note_dur = CYCLES_PER_US * 714;
		18: note_dur = CYCLES_PER_US * 342143;
		19: note_dur = CYCLES_PER_US * 714;
		20: note_dur = CYCLES_PER_US * 170714;
		21: note_dur = CYCLES_PER_US * 714;
		22: note_dur = CYCLES_PER_US * 170714;
		23: note_dur = CYCLES_PER_US * 714;
		24: note_dur = CYCLES_PER_US * 170714;
		25: note_dur = CYCLES_PER_US * 714;
		26: note_dur = CYCLES_PER_US * 170714;
		27: note_dur = CYCLES_PER_US * 172143;
		28: note_dur = CYCLES_PER_US * 170714;
		29: note_dur = CYCLES_PER_US * 1200714;
		30: note_dur = CYCLES_PER_US * 170714;
		31: note_dur = CYCLES_PER_US * 714;
		32: note_dur = CYCLES_PER_US * 342143;
		33: note_dur = CYCLES_PER_US * 714;
		34: note_dur = CYCLES_PER_US * 170714;
		35: note_dur = CYCLES_PER_US * 714;
		36: note_dur = CYCLES_PER_US * 170714;
		37: note_dur = CYCLES_PER_US * 714;
		38: note_dur = CYCLES_PER_US * 170714;
		39: note_dur = CYCLES_PER_US * 714;
		40: note_dur = CYCLES_PER_US * 170714;
		41: note_dur = CYCLES_PER_US * 172143;
		42: note_dur = CYCLES_PER_US * 170714;
		43: note_dur = CYCLES_PER_US * 172143;
		44: note_dur = CYCLES_PER_US * 170714;
		45: note_dur = CYCLES_PER_US * 857857;
		46: note_dur = CYCLES_PER_US * 170714;
		47: note_dur = CYCLES_PER_US * 714;
		48: note_dur = CYCLES_PER_US * 342143;
		49: note_dur = CYCLES_PER_US * 714;
		50: note_dur = CYCLES_PER_US * 170714;
		51: note_dur = CYCLES_PER_US * 714;
		52: note_dur = CYCLES_PER_US * 170714;
		53: note_dur = CYCLES_PER_US * 714;
		54: note_dur = CYCLES_PER_US * 170714;
		55: note_dur = CYCLES_PER_US * 714;
		56: note_dur = CYCLES_PER_US * 170714;
		57: note_dur = CYCLES_PER_US * 172143;
		58: note_dur = CYCLES_PER_US * 170714;
		59: note_dur = CYCLES_PER_US * 1372142;
		60: note_dur = CYCLES_PER_US * 342143;
		61: note_dur = CYCLES_PER_US * 714;
		62: note_dur = CYCLES_PER_US * 342143;
		63: note_dur = CYCLES_PER_US * 714;
		64: note_dur = CYCLES_PER_US * 427857;
		65: note_dur = CYCLES_PER_US * 714;
		66: note_dur = CYCLES_PER_US * 170714;
		67: note_dur = CYCLES_PER_US * 172143;
		68: note_dur = CYCLES_PER_US * 170714;
		69: note_dur = CYCLES_PER_US * 172143;
		70: note_dur = CYCLES_PER_US * 170714;
		71: note_dur = CYCLES_PER_US * 714;
		72: note_dur = CYCLES_PER_US * 170714;
		73: note_dur = CYCLES_PER_US * 714;
		74: note_dur = CYCLES_PER_US * 170714;
		75: note_dur = CYCLES_PER_US * 714;
		76: note_dur = CYCLES_PER_US * 342143;
		77: note_dur = CYCLES_PER_US * 714;
		78: note_dur = CYCLES_PER_US * 342143;
		79: note_dur = CYCLES_PER_US * 714;
		80: note_dur = CYCLES_PER_US * 342143;
		81: note_dur = CYCLES_PER_US * 714;
		82: note_dur = CYCLES_PER_US * 427857;
		83: note_dur = CYCLES_PER_US * 714;
		84: note_dur = CYCLES_PER_US * 170714;
		85: note_dur = CYCLES_PER_US * 172143;
		86: note_dur = CYCLES_PER_US * 170714;
		87: note_dur = CYCLES_PER_US * 172143;
		88: note_dur = CYCLES_PER_US * 170714;
		89: note_dur = CYCLES_PER_US * 714;
		90: note_dur = CYCLES_PER_US * 170714;
		91: note_dur = CYCLES_PER_US * 714;
		92: note_dur = CYCLES_PER_US * 170714;
		93: note_dur = CYCLES_PER_US * 714;
		94: note_dur = CYCLES_PER_US * 170714;
		95: note_dur = CYCLES_PER_US * 714;
		96: note_dur = CYCLES_PER_US * 170714;
		97: note_dur = CYCLES_PER_US * 714;
		98: note_dur = CYCLES_PER_US * 342143;
		99: note_dur = CYCLES_PER_US * 714;
		100: note_dur = CYCLES_PER_US * 342143;
		101: note_dur = CYCLES_PER_US * 714;
		102: note_dur = CYCLES_PER_US * 427857;
		103: note_dur = CYCLES_PER_US * 714;
		104: note_dur = CYCLES_PER_US * 170714;
		105: note_dur = CYCLES_PER_US * 172143;
		106: note_dur = CYCLES_PER_US * 170714;
		107: note_dur = CYCLES_PER_US * 172143;
		108: note_dur = CYCLES_PER_US * 170714;
		109: note_dur = CYCLES_PER_US * 714;
		110: note_dur = CYCLES_PER_US * 170714;
		111: note_dur = CYCLES_PER_US * 714;
		112: note_dur = CYCLES_PER_US * 170714;
		113: note_dur = CYCLES_PER_US * 714;
		114: note_dur = CYCLES_PER_US * 342143;
		115: note_dur = CYCLES_PER_US * 714;
		116: note_dur = CYCLES_PER_US * 342143;
		117: note_dur = CYCLES_PER_US * 714;
		118: note_dur = CYCLES_PER_US * 342143;
		119: note_dur = CYCLES_PER_US * 714;
		120: note_dur = CYCLES_PER_US * 427857;
		121: note_dur = CYCLES_PER_US * 714;
		122: note_dur = CYCLES_PER_US * 170714;
		123: note_dur = CYCLES_PER_US * 172143;
		124: note_dur = CYCLES_PER_US * 170714;
		125: note_dur = CYCLES_PER_US * 172143;
		126: note_dur = CYCLES_PER_US * 170714;
		127: note_dur = CYCLES_PER_US * 172143;
		128: note_dur = CYCLES_PER_US * 170714;
		129: note_dur = CYCLES_PER_US * 714;
		130: note_dur = CYCLES_PER_US * 170714;
		131: note_dur = CYCLES_PER_US * 714;
		132: note_dur = CYCLES_PER_US * 170714;
		133: note_dur = CYCLES_PER_US * 714;
		134: note_dur = CYCLES_PER_US * 1370714;
		135: note_dur = CYCLES_PER_US * 714;
		136: note_dur = CYCLES_PER_US * 342143;
		137: note_dur = CYCLES_PER_US * 172143;
		138: note_dur = CYCLES_PER_US * 85000;
		139: note_dur = CYCLES_PER_US * 172143;
		140: note_dur = CYCLES_PER_US * 170714;
		141: note_dur = CYCLES_PER_US * 714;
		142: note_dur = CYCLES_PER_US * 170714;
		143: note_dur = CYCLES_PER_US * 714;
		144: note_dur = CYCLES_PER_US * 170714;
		145: note_dur = CYCLES_PER_US * 714;
		146: note_dur = CYCLES_PER_US * 1370714;
		147: note_dur = CYCLES_PER_US * 714;
		148: note_dur = CYCLES_PER_US * 342143;
		149: note_dur = CYCLES_PER_US * 172143;
		150: note_dur = CYCLES_PER_US * 85000;
		151: note_dur = CYCLES_PER_US * 172143;
		152: note_dur = CYCLES_PER_US * 170714;
		153: note_dur = CYCLES_PER_US * 714;
		154: note_dur = CYCLES_PER_US * 170714;
		155: note_dur = CYCLES_PER_US * 714;
		156: note_dur = CYCLES_PER_US * 170714;
		157: note_dur = CYCLES_PER_US * 714;
		158: note_dur = CYCLES_PER_US * 1370714;
		159: note_dur = CYCLES_PER_US * 714;
		160: note_dur = CYCLES_PER_US * 342143;
		161: note_dur = CYCLES_PER_US * 172143;
		162: note_dur = CYCLES_PER_US * 85000;
		163: note_dur = CYCLES_PER_US * 686428;
		164: note_dur = CYCLES_PER_US * 170714;
		165: note_dur = CYCLES_PER_US * 714;
		166: note_dur = CYCLES_PER_US * 170714;
		167: note_dur = CYCLES_PER_US * 714;
		168: note_dur = CYCLES_PER_US * 170714;
		169: note_dur = CYCLES_PER_US * 714;
		170: note_dur = CYCLES_PER_US * 170714;
		171: note_dur = CYCLES_PER_US * 714;
		172: note_dur = CYCLES_PER_US * 342143;
		173: note_dur = CYCLES_PER_US * 714;
		174: note_dur = CYCLES_PER_US * 342143;
		175: note_dur = CYCLES_PER_US * 714;
		176: note_dur = CYCLES_PER_US * 256428;
		177: note_dur = CYCLES_PER_US * 514286;
		178: note_dur = CYCLES_PER_US * 342143;
		179: note_dur = CYCLES_PER_US * 714;
		180: note_dur = CYCLES_PER_US * 342143;
		181: note_dur = CYCLES_PER_US * 714;
		182: note_dur = CYCLES_PER_US * 427857;
		183: note_dur = CYCLES_PER_US * 714;
		184: note_dur = CYCLES_PER_US * 170714;
		185: note_dur = CYCLES_PER_US * 172143;
		186: note_dur = CYCLES_PER_US * 170714;
		187: note_dur = CYCLES_PER_US * 172143;
		188: note_dur = CYCLES_PER_US * 170714;
		189: note_dur = CYCLES_PER_US * 714;
		190: note_dur = CYCLES_PER_US * 170714;
		191: note_dur = CYCLES_PER_US * 714;
		192: note_dur = CYCLES_PER_US * 170714;
		193: note_dur = CYCLES_PER_US * 714;
		194: note_dur = CYCLES_PER_US * 342143;
		195: note_dur = CYCLES_PER_US * 714;
		196: note_dur = CYCLES_PER_US * 342143;
		197: note_dur = CYCLES_PER_US * 714;
		198: note_dur = CYCLES_PER_US * 342143;
		199: note_dur = CYCLES_PER_US * 714;
		200: note_dur = CYCLES_PER_US * 427857;
		201: note_dur = CYCLES_PER_US * 714;
		202: note_dur = CYCLES_PER_US * 170714;
		203: note_dur = CYCLES_PER_US * 172143;
		204: note_dur = CYCLES_PER_US * 170714;
		205: note_dur = CYCLES_PER_US * 172143;
		206: note_dur = CYCLES_PER_US * 170714;
		207: note_dur = CYCLES_PER_US * 714;
		208: note_dur = CYCLES_PER_US * 170714;
		209: note_dur = CYCLES_PER_US * 714;
		210: note_dur = CYCLES_PER_US * 170714;
		211: note_dur = CYCLES_PER_US * 714;
		212: note_dur = CYCLES_PER_US * 170714;
		213: note_dur = CYCLES_PER_US * 714;
		214: note_dur = CYCLES_PER_US * 170714;
		215: note_dur = CYCLES_PER_US * 714;
		216: note_dur = CYCLES_PER_US * 342143;
		217: note_dur = CYCLES_PER_US * 714;
		218: note_dur = CYCLES_PER_US * 342143;
		219: note_dur = CYCLES_PER_US * 714;
		220: note_dur = CYCLES_PER_US * 427857;
		221: note_dur = CYCLES_PER_US * 714;
		222: note_dur = CYCLES_PER_US * 170714;
		223: note_dur = CYCLES_PER_US * 172143;
		224: note_dur = CYCLES_PER_US * 170714;
		225: note_dur = CYCLES_PER_US * 172143;
		226: note_dur = CYCLES_PER_US * 170714;
		227: note_dur = CYCLES_PER_US * 714;
		228: note_dur = CYCLES_PER_US * 170714;
		229: note_dur = CYCLES_PER_US * 714;
		230: note_dur = CYCLES_PER_US * 170714;
		231: note_dur = CYCLES_PER_US * 714;
		232: note_dur = CYCLES_PER_US * 342143;
		233: note_dur = CYCLES_PER_US * 714;
		234: note_dur = CYCLES_PER_US * 342143;
		235: note_dur = CYCLES_PER_US * 714;
		236: note_dur = CYCLES_PER_US * 342143;
		237: note_dur = CYCLES_PER_US * 714;
		238: note_dur = CYCLES_PER_US * 427857;
		239: note_dur = CYCLES_PER_US * 714;
		240: note_dur = CYCLES_PER_US * 170714;
		241: note_dur = CYCLES_PER_US * 915000;
		242: note_dur = CYCLES_PER_US * 227857;
		243: note_dur = CYCLES_PER_US * 714;
		244: note_dur = CYCLES_PER_US * 227857;
		245: note_dur = CYCLES_PER_US * 714;
		246: note_dur = CYCLES_PER_US * 227857;
		247: note_dur = CYCLES_PER_US * 714;
		248: note_dur = CYCLES_PER_US * 227857;
		249: note_dur = CYCLES_PER_US * 714;
		250: note_dur = CYCLES_PER_US * 227857;
		251: note_dur = CYCLES_PER_US * 714;
		252: note_dur = CYCLES_PER_US * 170714;
		253: note_dur = CYCLES_PER_US * 714;
		254: note_dur = CYCLES_PER_US * 170714;
		255: note_dur = CYCLES_PER_US * 714;
		256: note_dur = CYCLES_PER_US * 170714;
		257: note_dur = CYCLES_PER_US * 714;
		258: note_dur = CYCLES_PER_US * 342143;
		259: note_dur = CYCLES_PER_US * 714;
		260: note_dur = CYCLES_PER_US * 742143;
		261: note_dur = CYCLES_PER_US * 714;
		262: note_dur = CYCLES_PER_US * 227857;
		263: note_dur = CYCLES_PER_US * 714;
		264: note_dur = CYCLES_PER_US * 227857;
		265: note_dur = CYCLES_PER_US * 714;
		266: note_dur = CYCLES_PER_US * 227857;
		267: note_dur = CYCLES_PER_US * 714;
		268: note_dur = CYCLES_PER_US * 227857;
		269: note_dur = CYCLES_PER_US * 714;
		270: note_dur = CYCLES_PER_US * 227857;
		271: note_dur = CYCLES_PER_US * 714;
		272: note_dur = CYCLES_PER_US * 170714;
		273: note_dur = CYCLES_PER_US * 714;
		274: note_dur = CYCLES_PER_US * 85000;
		275: note_dur = CYCLES_PER_US * 714;
		276: note_dur = CYCLES_PER_US * 85000;
		277: note_dur = CYCLES_PER_US * 714;
		278: note_dur = CYCLES_PER_US * 170714;
		279: note_dur = CYCLES_PER_US * 714;
		280: note_dur = CYCLES_PER_US * 513571;
		281: note_dur = CYCLES_PER_US * 857857;
		282: note_dur = CYCLES_PER_US * 170714;
		283: note_dur = CYCLES_PER_US * 714;
		284: note_dur = CYCLES_PER_US * 170714;
		285: note_dur = CYCLES_PER_US * 714;
		286: note_dur = CYCLES_PER_US * 170714;
		287: note_dur = CYCLES_PER_US * 714;
		288: note_dur = CYCLES_PER_US * 714;
		289: note_dur = CYCLES_PER_US * 0;
		290: note_dur = CYCLES_PER_US * 67857;
		291: note_dur = CYCLES_PER_US * 714;
		292: note_dur = CYCLES_PER_US * 67857;
		293: note_dur = CYCLES_PER_US * 714;
		294: note_dur = CYCLES_PER_US * 136429;
		295: note_dur = CYCLES_PER_US * 0;
		296: note_dur = CYCLES_PER_US * 714;
		297: note_dur = CYCLES_PER_US * 0;
		298: note_dur = CYCLES_PER_US * 85000;
		299: note_dur = CYCLES_PER_US * 714;
		300: note_dur = CYCLES_PER_US * 170714;
		301: note_dur = CYCLES_PER_US * 714;
		302: note_dur = CYCLES_PER_US * 714;
		303: note_dur = CYCLES_PER_US * 0;
		304: note_dur = CYCLES_PER_US * 67857;
		305: note_dur = CYCLES_PER_US * 714;
		306: note_dur = CYCLES_PER_US * 67857;
		307: note_dur = CYCLES_PER_US * 714;
		308: note_dur = CYCLES_PER_US * 136429;
		309: note_dur = CYCLES_PER_US * 714;
		310: note_dur = CYCLES_PER_US * 67857;
		311: note_dur = CYCLES_PER_US * 714;
		312: note_dur = CYCLES_PER_US * 67857;
		313: note_dur = CYCLES_PER_US * 714;
		314: note_dur = CYCLES_PER_US * 67857;
		315: note_dur = CYCLES_PER_US * 714;
		316: note_dur = CYCLES_PER_US * 136429;
		317: note_dur = CYCLES_PER_US * 714;
		318: note_dur = CYCLES_PER_US * 67857;
		319: note_dur = CYCLES_PER_US * 714;
		320: note_dur = CYCLES_PER_US * 67857;
		321: note_dur = CYCLES_PER_US * 714;
		322: note_dur = CYCLES_PER_US * 67857;
		323: note_dur = CYCLES_PER_US * 714;
		324: note_dur = CYCLES_PER_US * 136429;
		325: note_dur = CYCLES_PER_US * 714;
		326: note_dur = CYCLES_PER_US * 67857;
		327: note_dur = CYCLES_PER_US * 714;
		328: note_dur = CYCLES_PER_US * 67857;
		329: note_dur = CYCLES_PER_US * 714;
		330: note_dur = CYCLES_PER_US * 67857;
		331: note_dur = CYCLES_PER_US * 714;
		332: note_dur = CYCLES_PER_US * 136429;
		333: note_dur = CYCLES_PER_US * 714;
		334: note_dur = CYCLES_PER_US * 67857;
		335: note_dur = CYCLES_PER_US * 714;
		336: note_dur = CYCLES_PER_US * 67857;
		337: note_dur = CYCLES_PER_US * 714;
		338: note_dur = CYCLES_PER_US * 67857;
		339: note_dur = CYCLES_PER_US * 714;
		340: note_dur = CYCLES_PER_US * 136429;
		341: note_dur = CYCLES_PER_US * 0;
		342: note_dur = CYCLES_PER_US * 256428;
		343: note_dur = CYCLES_PER_US * 714;
		344: note_dur = CYCLES_PER_US * 170714;
		345: note_dur = CYCLES_PER_US * 714;
		346: note_dur = CYCLES_PER_US * 170714;
		347: note_dur = CYCLES_PER_US * 714;
		348: note_dur = CYCLES_PER_US * 170714;
		349: note_dur = CYCLES_PER_US * 714;
		350: note_dur = CYCLES_PER_US * 170714;
		351: note_dur = CYCLES_PER_US * 714;
		352: note_dur = CYCLES_PER_US * 170714;
		353: note_dur = CYCLES_PER_US * 714;
		354: note_dur = CYCLES_PER_US * 170714;
		355: note_dur = CYCLES_PER_US * 857857;
		356: note_dur = CYCLES_PER_US * 1713571;
		357: note_dur = CYCLES_PER_US * 714;
		358: note_dur = CYCLES_PER_US * 170714;
		359: note_dur = CYCLES_PER_US * 714;
		360: note_dur = CYCLES_PER_US * 85000;
		361: note_dur = CYCLES_PER_US * 714;
		362: note_dur = CYCLES_PER_US * 85000;
		363: note_dur = CYCLES_PER_US * 714;
		364: note_dur = CYCLES_PER_US * 85000;
		365: note_dur = CYCLES_PER_US * 714;
		366: note_dur = CYCLES_PER_US * 85000;
		367: note_dur = CYCLES_PER_US * 714;
		368: note_dur = CYCLES_PER_US * 85000;
		369: note_dur = CYCLES_PER_US * 714;
		370: note_dur = CYCLES_PER_US * 85000;
		371: note_dur = CYCLES_PER_US * 714;
		372: note_dur = CYCLES_PER_US * 85000;
		373: note_dur = CYCLES_PER_US * 714;
		374: note_dur = CYCLES_PER_US * 85000;
		375: note_dur = CYCLES_PER_US * 714;
		376: note_dur = CYCLES_PER_US * 85000;
		377: note_dur = CYCLES_PER_US * 714;
		378: note_dur = CYCLES_PER_US * 85000;
		379: note_dur = CYCLES_PER_US * 714;
		380: note_dur = CYCLES_PER_US * 85000;
		381: note_dur = CYCLES_PER_US * 714;
		382: note_dur = CYCLES_PER_US * 85000;
		383: note_dur = CYCLES_PER_US * 714;
		384: note_dur = CYCLES_PER_US * 85000;
		385: note_dur = CYCLES_PER_US * 714;
		386: note_dur = CYCLES_PER_US * 85000;
		387: note_dur = CYCLES_PER_US * 714;
		388: note_dur = CYCLES_PER_US * 85000;
		389: note_dur = CYCLES_PER_US * 714;
		390: note_dur = CYCLES_PER_US * 85000;
		391: note_dur = CYCLES_PER_US * 714;
		392: note_dur = CYCLES_PER_US * 1199285;
		393: note_dur = CYCLES_PER_US * 714;
		394: note_dur = CYCLES_PER_US * 170714;
		395: note_dur = CYCLES_PER_US * 857857;
		396: note_dur = CYCLES_PER_US * 170714;
		397: note_dur = CYCLES_PER_US * 714;
		398: note_dur = CYCLES_PER_US * 570714;
		399: note_dur = CYCLES_PER_US * 714;
		400: note_dur = CYCLES_PER_US * 227857;
		401: note_dur = CYCLES_PER_US * 714;
		402: note_dur = CYCLES_PER_US * 227857;
		403: note_dur = CYCLES_PER_US * 714;
		404: note_dur = CYCLES_PER_US * 227857;
		405: note_dur = CYCLES_PER_US * 714;
		406: note_dur = CYCLES_PER_US * 227857;
		407: note_dur = CYCLES_PER_US * 714;
		408: note_dur = CYCLES_PER_US * 227857;
		409: note_dur = CYCLES_PER_US * 714;
		410: note_dur = CYCLES_PER_US * 227857;
		411: note_dur = CYCLES_PER_US * 714;
		412: note_dur = CYCLES_PER_US * 227857;
		413: note_dur = CYCLES_PER_US * 714;
		414: note_dur = CYCLES_PER_US * 227857;
		415: note_dur = CYCLES_PER_US * 714;
		416: note_dur = CYCLES_PER_US * 170714;
		417: note_dur = CYCLES_PER_US * 714;
		418: note_dur = CYCLES_PER_US * 85000;
		419: note_dur = CYCLES_PER_US * 714;
		420: note_dur = CYCLES_PER_US * 85000;
		421: note_dur = CYCLES_PER_US * 714;
		422: note_dur = CYCLES_PER_US * 170714;
		423: note_dur = CYCLES_PER_US * 714;
		424: note_dur = CYCLES_PER_US * 170714;
		425: note_dur = CYCLES_PER_US * 714;
		426: note_dur = CYCLES_PER_US * 342143;
		427: note_dur = CYCLES_PER_US * 714;
		428: note_dur = CYCLES_PER_US * 170714;
		429: note_dur = CYCLES_PER_US * 714;
		430: note_dur = CYCLES_PER_US * 85000;
		431: note_dur = CYCLES_PER_US * 714;
		432: note_dur = CYCLES_PER_US * 85000;
		433: note_dur = CYCLES_PER_US * 714;
		434: note_dur = CYCLES_PER_US * 170714;
		435: note_dur = CYCLES_PER_US * 714;
		436: note_dur = CYCLES_PER_US * 342143;
		437: note_dur = CYCLES_PER_US * 714;
		438: note_dur = CYCLES_PER_US * 513571;
		439: note_dur = CYCLES_PER_US * 515000;
		440: note_dur = CYCLES_PER_US * 170714;
		441: note_dur = CYCLES_PER_US * 714;
		442: note_dur = CYCLES_PER_US * 170714;
		443: note_dur = CYCLES_PER_US * 714;
		444: note_dur = CYCLES_PER_US * 170714;
		445: note_dur = CYCLES_PER_US * 714;
		446: note_dur = CYCLES_PER_US * 1370714;
		447: note_dur = CYCLES_PER_US * 714;
		448: note_dur = CYCLES_PER_US * 342143;
		449: note_dur = CYCLES_PER_US * 172143;
		450: note_dur = CYCLES_PER_US * 85000;
		451: note_dur = CYCLES_PER_US * 172143;
		452: note_dur = CYCLES_PER_US * 170714;
		453: note_dur = CYCLES_PER_US * 714;
		454: note_dur = CYCLES_PER_US * 170714;
		455: note_dur = CYCLES_PER_US * 714;
		456: note_dur = CYCLES_PER_US * 170714;
		457: note_dur = CYCLES_PER_US * 714;
		458: note_dur = CYCLES_PER_US * 1370714;
		459: note_dur = CYCLES_PER_US * 714;
		460: note_dur = CYCLES_PER_US * 342143;
		461: note_dur = CYCLES_PER_US * 172143;
		462: note_dur = CYCLES_PER_US * 85000;
		463: note_dur = CYCLES_PER_US * 172143;
		464: note_dur = CYCLES_PER_US * 170714;
		465: note_dur = CYCLES_PER_US * 714;
		466: note_dur = CYCLES_PER_US * 170714;
		467: note_dur = CYCLES_PER_US * 714;
		468: note_dur = CYCLES_PER_US * 170714;
		469: note_dur = CYCLES_PER_US * 714;
		470: note_dur = CYCLES_PER_US * 1370714;
		471: note_dur = CYCLES_PER_US * 714;
		472: note_dur = CYCLES_PER_US * 342143;
		473: note_dur = CYCLES_PER_US * 172143;
		474: note_dur = CYCLES_PER_US * 85000;
		475: note_dur = CYCLES_PER_US * 686428;
		476: note_dur = CYCLES_PER_US * 170714;
		477: note_dur = CYCLES_PER_US * 714;
		478: note_dur = CYCLES_PER_US * 170714;
		479: note_dur = CYCLES_PER_US * 714;
		480: note_dur = CYCLES_PER_US * 170714;
		481: note_dur = CYCLES_PER_US * 714;
		482: note_dur = CYCLES_PER_US * 170714;
		483: note_dur = CYCLES_PER_US * 714;
		484: note_dur = CYCLES_PER_US * 342143;
		485: note_dur = CYCLES_PER_US * 714;
		486: note_dur = CYCLES_PER_US * 342143;
		487: note_dur = CYCLES_PER_US * 714;
		488: note_dur = CYCLES_PER_US * 256428;
		489: note_dur = CYCLES_PER_US * 342857;
		490: note_dur = CYCLES_PER_US * 170714;
		491: note_dur = CYCLES_PER_US * 714;
		492: note_dur = CYCLES_PER_US * 342143;
		493: note_dur = CYCLES_PER_US * 714;
		494: note_dur = CYCLES_PER_US * 170714;
		495: note_dur = CYCLES_PER_US * 714;
		496: note_dur = CYCLES_PER_US * 170714;
		497: note_dur = CYCLES_PER_US * 714;
		498: note_dur = CYCLES_PER_US * 170714;
		499: note_dur = CYCLES_PER_US * 172143;
		500: note_dur = CYCLES_PER_US * 170714;
		501: note_dur = CYCLES_PER_US * 714;
		502: note_dur = CYCLES_PER_US * 170714;
		503: note_dur = CYCLES_PER_US * 172143;
		504: note_dur = CYCLES_PER_US * 170714;
		505: note_dur = CYCLES_PER_US * 857857;
		506: note_dur = CYCLES_PER_US * 170714;
		507: note_dur = CYCLES_PER_US * 714;
		508: note_dur = CYCLES_PER_US * 342143;
		509: note_dur = CYCLES_PER_US * 714;
		510: note_dur = CYCLES_PER_US * 170714;
		511: note_dur = CYCLES_PER_US * 714;
		512: note_dur = CYCLES_PER_US * 170714;
		513: note_dur = CYCLES_PER_US * 714;
		514: note_dur = CYCLES_PER_US * 170714;
		515: note_dur = CYCLES_PER_US * 714;
		516: note_dur = CYCLES_PER_US * 170714;
		517: note_dur = CYCLES_PER_US * 172143;
		518: note_dur = CYCLES_PER_US * 170714;
		519: note_dur = CYCLES_PER_US * 1200714;
		520: note_dur = CYCLES_PER_US * 170714;
		521: note_dur = CYCLES_PER_US * 714;
		522: note_dur = CYCLES_PER_US * 342143;
		523: note_dur = CYCLES_PER_US * 714;
		524: note_dur = CYCLES_PER_US * 170714;
		525: note_dur = CYCLES_PER_US * 714;
		526: note_dur = CYCLES_PER_US * 170714;
		527: note_dur = CYCLES_PER_US * 714;
		528: note_dur = CYCLES_PER_US * 170714;
		529: note_dur = CYCLES_PER_US * 714;
		530: note_dur = CYCLES_PER_US * 170714;
		531: note_dur = CYCLES_PER_US * 172143;
		532: note_dur = CYCLES_PER_US * 170714;
		533: note_dur = CYCLES_PER_US * 172143;
		534: note_dur = CYCLES_PER_US * 170714;
		535: note_dur = CYCLES_PER_US * 857857;
		536: note_dur = CYCLES_PER_US * 170714;
		537: note_dur = CYCLES_PER_US * 714;
		538: note_dur = CYCLES_PER_US * 342143;
		539: note_dur = CYCLES_PER_US * 714;
		540: note_dur = CYCLES_PER_US * 170714;
		541: note_dur = CYCLES_PER_US * 714;
		542: note_dur = CYCLES_PER_US * 170714;
		543: note_dur = CYCLES_PER_US * 714;
		544: note_dur = CYCLES_PER_US * 170714;
		545: note_dur = CYCLES_PER_US * 714;
		546: note_dur = CYCLES_PER_US * 170714;
		547: note_dur = CYCLES_PER_US * 172143;
		548: note_dur = CYCLES_PER_US * 170714;
		549: note_dur = CYCLES_PER_US * 342857;
		550: note_dur = CYCLES_PER_US * 342143;
		551: note_dur = CYCLES_PER_US * 714;
		552: note_dur = CYCLES_PER_US * 427857;
		553: note_dur = CYCLES_PER_US * 714;
		554: note_dur = CYCLES_PER_US * 170714;
		555: note_dur = CYCLES_PER_US * 172143;
		556: note_dur = CYCLES_PER_US * 170714;
		557: note_dur = CYCLES_PER_US * 172143;
		558: note_dur = CYCLES_PER_US * 170714;
		559: note_dur = CYCLES_PER_US * 714;
		560: note_dur = CYCLES_PER_US * 170714;
		561: note_dur = CYCLES_PER_US * 714;
		562: note_dur = CYCLES_PER_US * 170714;
		563: note_dur = CYCLES_PER_US * 714;
		564: note_dur = CYCLES_PER_US * 342143;
		565: note_dur = CYCLES_PER_US * 343571;
		566: note_dur = CYCLES_PER_US * 342143;
		567: note_dur = CYCLES_PER_US * 714;
		568: note_dur = CYCLES_PER_US * 427857;
		569: note_dur = CYCLES_PER_US * 714;
		570: note_dur = CYCLES_PER_US * 170714;
		571: note_dur = CYCLES_PER_US * 172143;
		572: note_dur = CYCLES_PER_US * 170714;
		573: note_dur = CYCLES_PER_US * 172143;
		574: note_dur = CYCLES_PER_US * 170714;
		575: note_dur = CYCLES_PER_US * 714;
		576: note_dur = CYCLES_PER_US * 170714;
		577: note_dur = CYCLES_PER_US * 714;
		578: note_dur = CYCLES_PER_US * 170714;
		579: note_dur = CYCLES_PER_US * 714;
		580: note_dur = CYCLES_PER_US * 342143;
		581: note_dur = CYCLES_PER_US * 343571;
		582: note_dur = CYCLES_PER_US * 342143;
		583: note_dur = CYCLES_PER_US * 714;
		584: note_dur = CYCLES_PER_US * 427857;
		585: note_dur = CYCLES_PER_US * 714;
		586: note_dur = CYCLES_PER_US * 170714;
		587: note_dur = CYCLES_PER_US * 172143;
		588: note_dur = CYCLES_PER_US * 170714;
		589: note_dur = CYCLES_PER_US * 172143;
		590: note_dur = CYCLES_PER_US * 170714;
		591: note_dur = CYCLES_PER_US * 714;
		592: note_dur = CYCLES_PER_US * 170714;
		593: note_dur = CYCLES_PER_US * 714;
		594: note_dur = CYCLES_PER_US * 170714;
		595: note_dur = CYCLES_PER_US * 714;
		596: note_dur = CYCLES_PER_US * 342143;
		597: note_dur = CYCLES_PER_US * 343571;
		598: note_dur = CYCLES_PER_US * 342143;
		599: note_dur = CYCLES_PER_US * 714;
		600: note_dur = CYCLES_PER_US * 427857;
		601: note_dur = CYCLES_PER_US * 714;
		602: note_dur = CYCLES_PER_US * 170714;
		603: note_dur = CYCLES_PER_US * 172143;
		604: note_dur = CYCLES_PER_US * 170714;
		605: note_dur = CYCLES_PER_US * 172143;
		606: note_dur = CYCLES_PER_US * 170714;
		607: note_dur = CYCLES_PER_US * 714;
		608: note_dur = CYCLES_PER_US * 170714;
		609: note_dur = CYCLES_PER_US * 714;
		610: note_dur = CYCLES_PER_US * 170714;
		611: note_dur = CYCLES_PER_US * 714;
		612: note_dur = CYCLES_PER_US * 342143;
		613: note_dur = CYCLES_PER_US * 343571;
		614: note_dur = CYCLES_PER_US * 342143;
		615: note_dur = CYCLES_PER_US * 714;
		616: note_dur = CYCLES_PER_US * 427857;
		617: note_dur = CYCLES_PER_US * 714;
		618: note_dur = CYCLES_PER_US * 170714;
		619: note_dur = CYCLES_PER_US * 172143;
		620: note_dur = CYCLES_PER_US * 170714;
		621: note_dur = CYCLES_PER_US * 172143;
		622: note_dur = CYCLES_PER_US * 170714;
		623: note_dur = CYCLES_PER_US * 714;
		624: note_dur = CYCLES_PER_US * 170714;
		625: note_dur = CYCLES_PER_US * 714;
		626: note_dur = CYCLES_PER_US * 170714;
		627: note_dur = CYCLES_PER_US * 714;
		628: note_dur = CYCLES_PER_US * 342143;
		629: note_dur = CYCLES_PER_US * 343571;
		630: note_dur = CYCLES_PER_US * 342143;
		631: note_dur = CYCLES_PER_US * 714;
		632: note_dur = CYCLES_PER_US * 427857;
		633: note_dur = CYCLES_PER_US * 714;
		634: note_dur = CYCLES_PER_US * 170714;
		635: note_dur = CYCLES_PER_US * 172143;
		636: note_dur = CYCLES_PER_US * 170714;
		637: note_dur = CYCLES_PER_US * 172143;
		638: note_dur = CYCLES_PER_US * 170714;
		639: note_dur = CYCLES_PER_US * 714;
		640: note_dur = CYCLES_PER_US * 170714;
		641: note_dur = CYCLES_PER_US * 714;
		642: note_dur = CYCLES_PER_US * 170714;
		643: note_dur = CYCLES_PER_US * 714;
		644: note_dur = CYCLES_PER_US * 342143;
		645: note_dur = CYCLES_PER_US * 343571;
		646: note_dur = CYCLES_PER_US * 342143;
		647: note_dur = CYCLES_PER_US * 714;
		648: note_dur = CYCLES_PER_US * 427857;
		649: note_dur = CYCLES_PER_US * 714;
		650: note_dur = CYCLES_PER_US * 170714;
		651: note_dur = CYCLES_PER_US * 172143;
		652: note_dur = CYCLES_PER_US * 170714;
		653: note_dur = CYCLES_PER_US * 172143;
		654: note_dur = CYCLES_PER_US * 170714;
		655: note_dur = CYCLES_PER_US * 714;
		656: note_dur = CYCLES_PER_US * 170714;
		657: note_dur = CYCLES_PER_US * 714;
		658: note_dur = CYCLES_PER_US * 170714;
		659: note_dur = CYCLES_PER_US * 714;
		660: note_dur = CYCLES_PER_US * 342143;
		661: note_dur = CYCLES_PER_US * 343571;
		662: note_dur = CYCLES_PER_US * 342143;
		663: note_dur = CYCLES_PER_US * 714;
		664: note_dur = CYCLES_PER_US * 427857;
		665: note_dur = CYCLES_PER_US * 714;
		666: note_dur = CYCLES_PER_US * 170714;
		667: note_dur = CYCLES_PER_US * 172143;
		668: note_dur = CYCLES_PER_US * 170714;
		669: note_dur = CYCLES_PER_US * 172143;
		670: note_dur = CYCLES_PER_US * 170714;
		671: note_dur = CYCLES_PER_US * 172143;
		672: note_dur = CYCLES_PER_US * 170714;
		673: note_dur = CYCLES_PER_US * 714;
		674: note_dur = CYCLES_PER_US * 170714;
		675: note_dur = CYCLES_PER_US * 714;
		676: note_dur = CYCLES_PER_US * 170714;
		677: note_dur = CYCLES_PER_US * 714;
		678: note_dur = CYCLES_PER_US * 1370714;
		679: note_dur = CYCLES_PER_US * 714;
		680: note_dur = CYCLES_PER_US * 342143;
		681: note_dur = CYCLES_PER_US * 172143;
		682: note_dur = CYCLES_PER_US * 85000;
		683: note_dur = CYCLES_PER_US * 172143;
		684: note_dur = CYCLES_PER_US * 170714;
		685: note_dur = CYCLES_PER_US * 714;
		686: note_dur = CYCLES_PER_US * 170714;
		687: note_dur = CYCLES_PER_US * 714;
		688: note_dur = CYCLES_PER_US * 170714;
		689: note_dur = CYCLES_PER_US * 714;
		690: note_dur = CYCLES_PER_US * 1370714;
		691: note_dur = CYCLES_PER_US * 714;
		692: note_dur = CYCLES_PER_US * 342143;
		693: note_dur = CYCLES_PER_US * 172143;
		694: note_dur = CYCLES_PER_US * 85000;
		695: note_dur = CYCLES_PER_US * 172143;
		696: note_dur = CYCLES_PER_US * 170714;
		697: note_dur = CYCLES_PER_US * 714;
		698: note_dur = CYCLES_PER_US * 170714;
		699: note_dur = CYCLES_PER_US * 714;
		700: note_dur = CYCLES_PER_US * 170714;
		701: note_dur = CYCLES_PER_US * 714;
		702: note_dur = CYCLES_PER_US * 1370714;
		703: note_dur = CYCLES_PER_US * 714;
		704: note_dur = CYCLES_PER_US * 342143;
		705: note_dur = CYCLES_PER_US * 172143;
		706: note_dur = CYCLES_PER_US * 85000;
		707: note_dur = CYCLES_PER_US * 686428;
		708: note_dur = CYCLES_PER_US * 170714;
		709: note_dur = CYCLES_PER_US * 714;
		710: note_dur = CYCLES_PER_US * 170714;
		711: note_dur = CYCLES_PER_US * 714;
		712: note_dur = CYCLES_PER_US * 170714;
		713: note_dur = CYCLES_PER_US * 714;
		714: note_dur = CYCLES_PER_US * 170714;
		715: note_dur = CYCLES_PER_US * 714;
		716: note_dur = CYCLES_PER_US * 342143;
		717: note_dur = CYCLES_PER_US * 714;
		718: note_dur = CYCLES_PER_US * 342143;
		719: note_dur = CYCLES_PER_US * 714;
		720: note_dur = CYCLES_PER_US * 256428;
		721: note_dur = CYCLES_PER_US * 342857;
		722: note_dur = CYCLES_PER_US * 170714;
		723: note_dur = CYCLES_PER_US * 714;
		724: note_dur = CYCLES_PER_US * 342143;
		725: note_dur = CYCLES_PER_US * 714;
		726: note_dur = CYCLES_PER_US * 170714;
		727: note_dur = CYCLES_PER_US * 714;
		728: note_dur = CYCLES_PER_US * 170714;
		729: note_dur = CYCLES_PER_US * 714;
		730: note_dur = CYCLES_PER_US * 170714;
		731: note_dur = CYCLES_PER_US * 172143;
		732: note_dur = CYCLES_PER_US * 170714;
		733: note_dur = CYCLES_PER_US * 714;
		734: note_dur = CYCLES_PER_US * 170714;
		735: note_dur = CYCLES_PER_US * 172143;
		736: note_dur = CYCLES_PER_US * 170714;
		737: note_dur = CYCLES_PER_US * 857857;
		738: note_dur = CYCLES_PER_US * 170714;
		739: note_dur = CYCLES_PER_US * 714;
		740: note_dur = CYCLES_PER_US * 342143;
		741: note_dur = CYCLES_PER_US * 714;
		742: note_dur = CYCLES_PER_US * 170714;
		743: note_dur = CYCLES_PER_US * 714;
		744: note_dur = CYCLES_PER_US * 170714;
		745: note_dur = CYCLES_PER_US * 714;
		746: note_dur = CYCLES_PER_US * 170714;
		747: note_dur = CYCLES_PER_US * 714;
		748: note_dur = CYCLES_PER_US * 170714;
		749: note_dur = CYCLES_PER_US * 172143;
		750: note_dur = CYCLES_PER_US * 170714;
		751: note_dur = CYCLES_PER_US * 1200714;
		752: note_dur = CYCLES_PER_US * 170714;
		753: note_dur = CYCLES_PER_US * 714;
		754: note_dur = CYCLES_PER_US * 342143;
		755: note_dur = CYCLES_PER_US * 714;
		756: note_dur = CYCLES_PER_US * 170714;
		757: note_dur = CYCLES_PER_US * 714;
		758: note_dur = CYCLES_PER_US * 170714;
		759: note_dur = CYCLES_PER_US * 714;
		760: note_dur = CYCLES_PER_US * 170714;
		761: note_dur = CYCLES_PER_US * 714;
		762: note_dur = CYCLES_PER_US * 170714;
		763: note_dur = CYCLES_PER_US * 172143;
		764: note_dur = CYCLES_PER_US * 170714;
		765: note_dur = CYCLES_PER_US * 172143;
		766: note_dur = CYCLES_PER_US * 170714;
		767: note_dur = CYCLES_PER_US * 857857;
		768: note_dur = CYCLES_PER_US * 170714;
		769: note_dur = CYCLES_PER_US * 714;
		770: note_dur = CYCLES_PER_US * 342143;
		771: note_dur = CYCLES_PER_US * 714;
		772: note_dur = CYCLES_PER_US * 170714;
		773: note_dur = CYCLES_PER_US * 714;
		774: note_dur = CYCLES_PER_US * 170714;
		775: note_dur = CYCLES_PER_US * 714;
		776: note_dur = CYCLES_PER_US * 170714;
		777: note_dur = CYCLES_PER_US * 714;
		778: note_dur = CYCLES_PER_US * 170714;
		779: note_dur = CYCLES_PER_US * 172143;
		780: note_dur = CYCLES_PER_US * 170714;
		781: note_dur = CYCLES_PER_US * 1372142;
		782: note_dur = CYCLES_PER_US * 342143;
		783: note_dur = CYCLES_PER_US * 714;
		784: note_dur = CYCLES_PER_US * 342143;
		785: note_dur = CYCLES_PER_US * 714;
		786: note_dur = CYCLES_PER_US * 427857;
		787: note_dur = CYCLES_PER_US * 714;
		788: note_dur = CYCLES_PER_US * 170714;
		789: note_dur = CYCLES_PER_US * 172143;
		790: note_dur = CYCLES_PER_US * 170714;
		791: note_dur = CYCLES_PER_US * 172143;
		792: note_dur = CYCLES_PER_US * 170714;
		793: note_dur = CYCLES_PER_US * 714;
		794: note_dur = CYCLES_PER_US * 170714;
		795: note_dur = CYCLES_PER_US * 714;
		796: note_dur = CYCLES_PER_US * 170714;
		797: note_dur = CYCLES_PER_US * 714;
		798: note_dur = CYCLES_PER_US * 342143;
		799: note_dur = CYCLES_PER_US * 714;
		800: note_dur = CYCLES_PER_US * 342143;
		801: note_dur = CYCLES_PER_US * 714;
		802: note_dur = CYCLES_PER_US * 342143;
		803: note_dur = CYCLES_PER_US * 714;
		804: note_dur = CYCLES_PER_US * 427857;
		805: note_dur = CYCLES_PER_US * 714;
		806: note_dur = CYCLES_PER_US * 170714;
		807: note_dur = CYCLES_PER_US * 172143;
		808: note_dur = CYCLES_PER_US * 170714;
		809: note_dur = CYCLES_PER_US * 172143;
		810: note_dur = CYCLES_PER_US * 170714;
		811: note_dur = CYCLES_PER_US * 714;
		812: note_dur = CYCLES_PER_US * 170714;
		813: note_dur = CYCLES_PER_US * 714;
		814: note_dur = CYCLES_PER_US * 170714;
		815: note_dur = CYCLES_PER_US * 714;
		816: note_dur = CYCLES_PER_US * 170714;
		817: note_dur = CYCLES_PER_US * 714;
		818: note_dur = CYCLES_PER_US * 170714;
		819: note_dur = CYCLES_PER_US * 714;
		820: note_dur = CYCLES_PER_US * 342143;
		821: note_dur = CYCLES_PER_US * 714;
		822: note_dur = CYCLES_PER_US * 342143;
		823: note_dur = CYCLES_PER_US * 714;
		824: note_dur = CYCLES_PER_US * 427857;
		825: note_dur = CYCLES_PER_US * 714;
		826: note_dur = CYCLES_PER_US * 170714;
		827: note_dur = CYCLES_PER_US * 172143;
		828: note_dur = CYCLES_PER_US * 170714;
		829: note_dur = CYCLES_PER_US * 172143;
		830: note_dur = CYCLES_PER_US * 170714;
		831: note_dur = CYCLES_PER_US * 714;
		832: note_dur = CYCLES_PER_US * 170714;
		833: note_dur = CYCLES_PER_US * 714;
		834: note_dur = CYCLES_PER_US * 170714;
		835: note_dur = CYCLES_PER_US * 714;
		836: note_dur = CYCLES_PER_US * 342143;
		837: note_dur = CYCLES_PER_US * 714;
		838: note_dur = CYCLES_PER_US * 342143;
		839: note_dur = CYCLES_PER_US * 714;
		840: note_dur = CYCLES_PER_US * 342143;
		841: note_dur = CYCLES_PER_US * 714;
		842: note_dur = CYCLES_PER_US * 427857;
		843: note_dur = CYCLES_PER_US * 714;
		844: note_dur = CYCLES_PER_US * 170714;
		845: note_dur = CYCLES_PER_US * 172143;
		846: note_dur = CYCLES_PER_US * 170714;
		847: note_dur = CYCLES_PER_US * 172143;
		848: note_dur = CYCLES_PER_US * 170714;
		849: note_dur = CYCLES_PER_US * 172143;
		850: note_dur = CYCLES_PER_US * 170714;
		851: note_dur = CYCLES_PER_US * 714;
		852: note_dur = CYCLES_PER_US * 170714;
		853: note_dur = CYCLES_PER_US * 714;
		854: note_dur = CYCLES_PER_US * 170714;
		855: note_dur = CYCLES_PER_US * 714;
		856: note_dur = CYCLES_PER_US * 1370714;
		857: note_dur = CYCLES_PER_US * 714;
		858: note_dur = CYCLES_PER_US * 342143;
		859: note_dur = CYCLES_PER_US * 172143;
		860: note_dur = CYCLES_PER_US * 85000;
		861: note_dur = CYCLES_PER_US * 172143;
		862: note_dur = CYCLES_PER_US * 170714;
		863: note_dur = CYCLES_PER_US * 714;
		864: note_dur = CYCLES_PER_US * 170714;
		865: note_dur = CYCLES_PER_US * 714;
		866: note_dur = CYCLES_PER_US * 170714;
		867: note_dur = CYCLES_PER_US * 714;
		868: note_dur = CYCLES_PER_US * 1370714;
		869: note_dur = CYCLES_PER_US * 714;
		870: note_dur = CYCLES_PER_US * 342143;
		871: note_dur = CYCLES_PER_US * 172143;
		872: note_dur = CYCLES_PER_US * 85000;
		873: note_dur = CYCLES_PER_US * 172143;
		874: note_dur = CYCLES_PER_US * 170714;
		875: note_dur = CYCLES_PER_US * 714;
		876: note_dur = CYCLES_PER_US * 170714;
		877: note_dur = CYCLES_PER_US * 714;
		878: note_dur = CYCLES_PER_US * 170714;
		879: note_dur = CYCLES_PER_US * 714;
		880: note_dur = CYCLES_PER_US * 1370714;
		881: note_dur = CYCLES_PER_US * 714;
		882: note_dur = CYCLES_PER_US * 342143;
		883: note_dur = CYCLES_PER_US * 172143;
		884: note_dur = CYCLES_PER_US * 85000;
		885: note_dur = CYCLES_PER_US * 686428;
		886: note_dur = CYCLES_PER_US * 170714;
		887: note_dur = CYCLES_PER_US * 714;
		888: note_dur = CYCLES_PER_US * 170714;
		889: note_dur = CYCLES_PER_US * 714;
		890: note_dur = CYCLES_PER_US * 170714;
		891: note_dur = CYCLES_PER_US * 714;
		892: note_dur = CYCLES_PER_US * 170714;
		893: note_dur = CYCLES_PER_US * 714;
		894: note_dur = CYCLES_PER_US * 342143;
		895: note_dur = CYCLES_PER_US * 714;
		896: note_dur = CYCLES_PER_US * 342143;
		897: note_dur = CYCLES_PER_US * 714;
		898: note_dur = CYCLES_PER_US * 256428;
		899: note_dur = CYCLES_PER_US * 342857;
		900: note_dur = CYCLES_PER_US * 170714;
		901: note_dur = CYCLES_PER_US * 714;
		902: note_dur = CYCLES_PER_US * 342143;
		903: note_dur = CYCLES_PER_US * 714;
		904: note_dur = CYCLES_PER_US * 342143;
		905: note_dur = CYCLES_PER_US * 714;
		906: note_dur = CYCLES_PER_US * 427857;
		907: note_dur = CYCLES_PER_US * 714;
		908: note_dur = CYCLES_PER_US * 170714;
		909: note_dur = CYCLES_PER_US * 172143;
		910: note_dur = CYCLES_PER_US * 170714;
		911: note_dur = CYCLES_PER_US * 172143;
		912: note_dur = CYCLES_PER_US * 170714;
		913: note_dur = CYCLES_PER_US * 714;
		914: note_dur = CYCLES_PER_US * 170714;
		915: note_dur = CYCLES_PER_US * 714;
		916: note_dur = CYCLES_PER_US * 170714;
		917: note_dur = CYCLES_PER_US * 714;
		918: note_dur = CYCLES_PER_US * 170714;
		919: note_dur = CYCLES_PER_US * 714;
		920: note_dur = CYCLES_PER_US * 170714;
		921: note_dur = CYCLES_PER_US * 714;
		922: note_dur = CYCLES_PER_US * 342143;
		923: note_dur = CYCLES_PER_US * 714;
		924: note_dur = CYCLES_PER_US * 170714;
		925: note_dur = CYCLES_PER_US * 714;
		926: note_dur = CYCLES_PER_US * 170714;
		927: note_dur = CYCLES_PER_US * 714;
		928: note_dur = CYCLES_PER_US * 170714;
		929: note_dur = CYCLES_PER_US * 714;
		930: note_dur = CYCLES_PER_US * 170714;
		931: note_dur = CYCLES_PER_US * 343571;
		932: note_dur = CYCLES_PER_US * 256428;
		933: note_dur = CYCLES_PER_US * 256428;
		default: note_dur = 0;
	endcase
end
endmodule